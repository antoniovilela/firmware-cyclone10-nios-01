// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition"

// DATE "09/17/2020 20:13:16"

// 
// Device: Altera 10CL016YU484C8G Package UFBGA484
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module processor (
	altera_reserved_tms,
	altera_reserved_tck,
	altera_reserved_tdi,
	altera_reserved_tdo,
	clk_clk,
	led_export,
	reset_reset_n,
	seg_export,
	seg_en_export,
	sw_export,
	uart_0_rxd,
	uart_0_txd)/* synthesis synthesis_greybox=1 */;
input 	altera_reserved_tms;
input 	altera_reserved_tck;
input 	altera_reserved_tdi;
output 	altera_reserved_tdo;
input 	clk_clk;
output 	[1:0] led_export;
input 	reset_reset_n;
output 	[7:0] seg_export;
output 	[2:0] seg_en_export;
input 	sw_export;
input 	uart_0_rxd;
output 	uart_0_txd;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[0]~q ;
wire \nios2_gen2_0|cpu|W_alu_result[7]~q ;
wire \nios2_gen2_0|cpu|W_alu_result[16]~q ;
wire \nios2_gen2_0|cpu|W_alu_result[15]~q ;
wire \nios2_gen2_0|cpu|W_alu_result[14]~q ;
wire \nios2_gen2_0|cpu|W_alu_result[13]~q ;
wire \nios2_gen2_0|cpu|W_alu_result[12]~q ;
wire \nios2_gen2_0|cpu|W_alu_result[11]~q ;
wire \nios2_gen2_0|cpu|W_alu_result[10]~q ;
wire \nios2_gen2_0|cpu|W_alu_result[9]~q ;
wire \nios2_gen2_0|cpu|W_alu_result[8]~q ;
wire \nios2_gen2_0|cpu|W_alu_result[4]~q ;
wire \nios2_gen2_0|cpu|W_alu_result[5]~q ;
wire \nios2_gen2_0|cpu|W_alu_result[6]~q ;
wire \nios2_gen2_0|cpu|W_alu_result[2]~q ;
wire \nios2_gen2_0|cpu|W_alu_result[3]~q ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[0] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[22] ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[22]~q ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[23] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[24] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[25] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[26] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[1] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[4] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[3] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[2] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[5] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[14] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[15] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[11] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[13] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[16] ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[16]~q ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[12] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[10] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[9] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[8] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[7] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[6] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[21] ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[21]~q ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[20] ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[20]~q ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[19] ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[19]~q ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[18] ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[18]~q ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[17] ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[17]~q ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[0]~q ;
wire \nios2_gen2_0|cpu|d_writedata[24]~q ;
wire \nios2_gen2_0|cpu|d_writedata[25]~q ;
wire \nios2_gen2_0|cpu|d_writedata[26]~q ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[1]~q ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[3]~q ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[2]~q ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[27] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[28] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[29] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[30] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[31] ;
wire \nios2_gen2_0|cpu|d_writedata[27]~q ;
wire \nios2_gen2_0|cpu|d_writedata[28]~q ;
wire \nios2_gen2_0|cpu|d_writedata[29]~q ;
wire \nios2_gen2_0|cpu|d_writedata[30]~q ;
wire \nios2_gen2_0|cpu|d_writedata[31]~q ;
wire \led|data_out[0]~q ;
wire \led|data_out[1]~q ;
wire \seg|data_out[0]~q ;
wire \seg|data_out[1]~q ;
wire \seg|data_out[2]~q ;
wire \seg|data_out[3]~q ;
wire \seg|data_out[4]~q ;
wire \seg|data_out[5]~q ;
wire \seg|data_out[6]~q ;
wire \seg|data_out[7]~q ;
wire \seg_en|data_out[0]~q ;
wire \seg_en|data_out[1]~q ;
wire \seg_en|data_out[2]~q ;
wire \uart_0|the_processor_uart_0_tx|txd~q ;
wire \jtag_uart_0|processor_jtag_uart_0_alt_jtag_atlantic|adapted_tdo~q ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_tck|ir_out[0]~q ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_tck|ir_out[1]~q ;
wire \nios2_gen2_0|cpu|d_writedata[0]~q ;
wire \rst_controller|r_sync_rst~q ;
wire \mm_interconnect_0|cmd_mux_003|saved_grant[0]~q ;
wire \nios2_gen2_0|cpu|d_write~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~0_combout ;
wire \mm_interconnect_0|cmd_mux_003|saved_grant[1]~q ;
wire \jtag_uart_0|processor_jtag_uart_0_alt_jtag_atlantic|rst1~q ;
wire \nios2_gen2_0|cpu|i_read~q ;
wire \nios2_gen2_0|cpu|F_pc[5]~q ;
wire \nios2_gen2_0|cpu|F_pc[14]~q ;
wire \nios2_gen2_0|cpu|F_pc[13]~q ;
wire \nios2_gen2_0|cpu|F_pc[12]~q ;
wire \nios2_gen2_0|cpu|F_pc[11]~q ;
wire \nios2_gen2_0|cpu|F_pc[10]~q ;
wire \nios2_gen2_0|cpu|F_pc[9]~q ;
wire \nios2_gen2_0|cpu|F_pc[8]~q ;
wire \nios2_gen2_0|cpu|F_pc[7]~q ;
wire \nios2_gen2_0|cpu|F_pc[6]~q ;
wire \nios2_gen2_0|cpu|F_pc[2]~q ;
wire \nios2_gen2_0|cpu|F_pc[3]~q ;
wire \nios2_gen2_0|cpu|F_pc[4]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_valid~3_combout ;
wire \nios2_gen2_0|cpu|d_read~q ;
wire \mm_interconnect_0|cmd_mux_003|src_valid~5_combout ;
wire \mm_interconnect_0|led_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \led|always0~0_combout ;
wire \nios2_gen2_0|cpu|F_pc[1]~q ;
wire \nios2_gen2_0|cpu|F_pc[0]~q ;
wire \sw|read_mux_out~0_combout ;
wire \sw|read_mux_out~1_combout ;
wire \mm_interconnect_0|led_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|led_s1_translator|wait_latency_counter[0]~q ;
wire \nios2_gen2_0|cpu|d_writedata[1]~q ;
wire \mm_interconnect_0|cmd_mux_005|saved_grant[0]~q ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~0_combout ;
wire \mm_interconnect_0|cmd_mux_005|saved_grant[1]~q ;
wire \mm_interconnect_0|cmd_mux_005|src_valid~2_combout ;
wire \mm_interconnect_0|cmd_mux_005|src_valid~4_combout ;
wire \mm_interconnect_0|seg_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \seg|always0~0_combout ;
wire \mm_interconnect_0|seg_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|seg_s1_translator|wait_latency_counter[0]~q ;
wire \nios2_gen2_0|cpu|d_writedata[2]~q ;
wire \nios2_gen2_0|cpu|d_writedata[3]~q ;
wire \nios2_gen2_0|cpu|d_writedata[4]~q ;
wire \nios2_gen2_0|cpu|d_writedata[5]~q ;
wire \nios2_gen2_0|cpu|d_writedata[6]~q ;
wire \nios2_gen2_0|cpu|d_writedata[7]~q ;
wire \mm_interconnect_0|cmd_mux_004|saved_grant[0]~q ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~0_combout ;
wire \mm_interconnect_0|cmd_mux_004|saved_grant[1]~q ;
wire \mm_interconnect_0|cmd_mux_004|src_valid~3_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_valid~5_combout ;
wire \mm_interconnect_0|seg_en_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \seg_en|always0~0_combout ;
wire \mm_interconnect_0|seg_en_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|seg_en_s1_translator|wait_latency_counter[0]~q ;
wire \mm_interconnect_0|rsp_demux|src0_valid~0_combout ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|read_latency_shift_reg[0]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|mem[0][74]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|mem[0][56]~q ;
wire \mm_interconnect_0|rsp_demux_001|src0_valid~0_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_translator|read_latency_shift_reg[0]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][74]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][56]~q ;
wire \mm_interconnect_0|rsp_demux_002|src0_valid~0_combout ;
wire \mm_interconnect_0|rsp_demux_003|src0_valid~0_combout ;
wire \mm_interconnect_0|rsp_mux|WideOr1~0_combout ;
wire \mm_interconnect_0|rsp_demux_004|src0_valid~0_combout ;
wire \mm_interconnect_0|seg_s1_translator|read_latency_shift_reg[0]~q ;
wire \mm_interconnect_0|seg_s1_agent_rsp_fifo|mem[0][74]~q ;
wire \mm_interconnect_0|seg_s1_agent_rsp_fifo|mem[0][56]~q ;
wire \mm_interconnect_0|rsp_demux_005|src0_valid~0_combout ;
wire \mm_interconnect_0|rsp_demux_007|src0_valid~0_combout ;
wire \mm_interconnect_0|rsp_mux|WideOr1~1_combout ;
wire \mm_interconnect_0|rsp_mux|WideOr1~combout ;
wire \mm_interconnect_0|cmd_mux_002|saved_grant[0]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|uart_0_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|uart_0_s1_translator|wait_latency_counter[1]~q ;
wire \jtag_uart_0|av_waitrequest~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|cmd_mux|saved_grant[0]~q ;
wire \mm_interconnect_0|cmd_mux_001|saved_grant[0]~q ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|the_processor_nios2_gen2_0_cpu_nios2_ocimem|waitrequest~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|cmd_mux_006|saved_grant[0]~q ;
wire \mm_interconnect_0|cmd_mux_006|saved_grant[1]~q ;
wire \mm_interconnect_0|nios2_gen2_0_data_master_translator|av_waitrequest~1_combout ;
wire \mm_interconnect_0|rsp_demux|src1_valid~0_combout ;
wire \mm_interconnect_0|rsp_demux_001|src1_valid~0_combout ;
wire \mm_interconnect_0|rsp_demux_002|src1_valid~0_combout ;
wire \mm_interconnect_0|rsp_demux_005|src1_valid~0_combout ;
wire \mm_interconnect_0|rsp_mux_001|WideOr1~0_combout ;
wire \mm_interconnect_0|rsp_demux_007|src1_valid~0_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~0_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~1_combout ;
wire \mm_interconnect_0|rsp_mux_001|WideOr1~1_combout ;
wire \mm_interconnect_0|nios2_gen2_0_data_master_translator|uav_write~0_combout ;
wire \nios2_gen2_0|cpu|d_writedata[9]~q ;
wire \mm_interconnect_0|cmd_mux_007|src_payload~0_combout ;
wire \mm_interconnect_0|cmd_mux_007|src_data[38]~combout ;
wire \mm_interconnect_0|cmd_mux_007|src_data[39]~combout ;
wire \mm_interconnect_0|cmd_mux_007|src_data[40]~combout ;
wire \mm_interconnect_0|cmd_mux_007|WideOr1~combout ;
wire \mm_interconnect_0|uart_0_s1_translator|av_begintransfer~0_combout ;
wire \mm_interconnect_0|cmd_mux|src_data[56]~combout ;
wire \mm_interconnect_0|cmd_mux|WideOr1~combout ;
wire \mm_interconnect_0|cmd_mux_001|WideOr1~combout ;
wire \mm_interconnect_0|cmd_mux_002|WideOr1~combout ;
wire \mm_interconnect_0|cmd_mux_007|src_data[56]~combout ;
wire \uart_0|the_processor_uart_0_rx|rx_rd_strobe_onset~0_combout ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_agent|rf_source_valid~0_combout ;
wire \nios2_gen2_0|cpu|hbreak_enabled~q ;
wire \mm_interconnect_0|rsp_mux|src_data[0]~combout ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[22]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[23]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[24]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[25]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[26]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_data[0]~0_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[0]~1_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[0]~3_combout ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[1]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[1]~q ;
wire \mm_interconnect_0|uart_0_s1_translator|av_readdata_pre[1]~q ;
wire \mm_interconnect_0|seg_s1_translator|av_readdata_pre[1]~q ;
wire \mm_interconnect_0|led_s1_translator|av_readdata_pre[1]~q ;
wire \mm_interconnect_0|seg_en_s1_translator|av_readdata_pre[1]~q ;
wire \mm_interconnect_0|seg_s1_translator|av_readdata_pre[4]~q ;
wire \mm_interconnect_0|uart_0_s1_translator|av_readdata_pre[4]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[4]~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[4]~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[3]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~4_combout ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[3]~q ;
wire \mm_interconnect_0|uart_0_s1_translator|av_readdata_pre[3]~q ;
wire \mm_interconnect_0|seg_s1_translator|av_readdata_pre[3]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[2]~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[2]~q ;
wire \mm_interconnect_0|seg_s1_translator|av_readdata_pre[2]~q ;
wire \mm_interconnect_0|seg_en_s1_translator|av_readdata_pre[2]~q ;
wire \mm_interconnect_0|uart_0_s1_translator|av_readdata_pre[2]~q ;
wire \mm_interconnect_0|cmd_mux_001|src_data[46]~combout ;
wire \mm_interconnect_0|seg_s1_translator|av_readdata_pre[5]~q ;
wire \mm_interconnect_0|uart_0_s1_translator|av_readdata_pre[5]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[5]~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[5]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[14]~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[14]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[15]~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[15]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~5_combout ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[11]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[13]~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[13]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[16]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[12]~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[12]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[10]~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[10]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[9]~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[9]~q ;
wire \mm_interconnect_0|uart_0_s1_translator|av_readdata_pre[9]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[8]~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[8]~q ;
wire \mm_interconnect_0|uart_0_s1_translator|av_readdata_pre[8]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[7]~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[7]~q ;
wire \mm_interconnect_0|seg_s1_translator|av_readdata_pre[7]~q ;
wire \mm_interconnect_0|uart_0_s1_translator|av_readdata_pre[7]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[6]~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[6]~q ;
wire \mm_interconnect_0|seg_s1_translator|av_readdata_pre[6]~q ;
wire \mm_interconnect_0|uart_0_s1_translator|av_readdata_pre[6]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[21]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[20]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[19]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[18]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[17]~q ;
wire \mm_interconnect_0|cmd_mux_007|src_payload~1_combout ;
wire \mm_interconnect_0|cmd_mux_007|src_payload~2_combout ;
wire \mm_interconnect_0|cmd_mux_007|src_payload~3_combout ;
wire \mm_interconnect_0|cmd_mux_007|src_payload~4_combout ;
wire \mm_interconnect_0|cmd_mux_007|src_payload~5_combout ;
wire \mm_interconnect_0|cmd_mux_007|src_payload~6_combout ;
wire \mm_interconnect_0|cmd_mux_007|src_payload~7_combout ;
wire \mm_interconnect_0|cmd_mux_007|src_payload~8_combout ;
wire \jtag_uart_0|the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_full~q ;
wire \rst_controller|r_early_rst~q ;
wire \mm_interconnect_0|rsp_mux|src_data[8]~5_combout ;
wire \seg|readdata[0]~combout ;
wire \seg_en|readdata[0]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~0_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[38]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[39]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[40]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[41]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[42]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[43]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[44]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[45]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[46]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[47]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[48]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[49]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[50]~combout ;
wire \nios2_gen2_0|cpu|d_byteenable[0]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_data[32]~combout ;
wire \jtag_uart_0|read_0~q ;
wire \jtag_uart_0|av_readdata[0]~0_combout ;
wire \uart_0|the_processor_uart_0_regs|readdata[0]~q ;
wire \led|readdata[0]~combout ;
wire \sw|readdata[0]~q ;
wire \jtag_uart_0|av_readdata[9]~combout ;
wire \jtag_uart_0|av_readdata[8]~1_combout ;
wire \uart_0|the_processor_uart_0_regs|irq~q ;
wire \nios2_gen2_0|cpu|d_writedata[22]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~1_combout ;
wire \nios2_gen2_0|cpu|d_byteenable[2]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_data[34]~combout ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[22]~q ;
wire \jtag_uart_0|the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_full~q ;
wire \jtag_uart_0|the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ;
wire \jtag_uart_0|the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ;
wire \jtag_uart_0|the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ;
wire \jtag_uart_0|the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ;
wire \jtag_uart_0|the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ;
wire \jtag_uart_0|the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[23]~q ;
wire \nios2_gen2_0|cpu|d_writedata[23]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~2_combout ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[24]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~3_combout ;
wire \nios2_gen2_0|cpu|d_byteenable[3]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_data[35]~combout ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[25]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~4_combout ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[26]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~5_combout ;
wire \jtag_uart_0|av_readdata[1]~2_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~6_combout ;
wire \uart_0|the_processor_uart_0_regs|readdata[1]~q ;
wire \seg|readdata[1]~combout ;
wire \led|readdata[1]~combout ;
wire \seg_en|readdata[1]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~7_combout ;
wire \seg|readdata[4]~combout ;
wire \uart_0|the_processor_uart_0_regs|readdata[4]~q ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[4]~q ;
wire \jtag_uart_0|av_readdata[4]~3_combout ;
wire \jtag_uart_0|av_readdata[3]~4_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~8_combout ;
wire \uart_0|the_processor_uart_0_regs|readdata[3]~q ;
wire \seg|readdata[3]~combout ;
wire \jtag_uart_0|av_readdata[2]~5_combout ;
wire \seg|readdata[2]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~9_combout ;
wire \seg_en|readdata[2]~combout ;
wire \uart_0|the_processor_uart_0_regs|readdata[2]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~10_combout ;
wire \seg|readdata[5]~combout ;
wire \uart_0|the_processor_uart_0_regs|readdata[5]~q ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[5]~q ;
wire \jtag_uart_0|av_readdata[5]~6_combout ;
wire \nios2_gen2_0|cpu|d_writedata[14]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~11_combout ;
wire \nios2_gen2_0|cpu|d_byteenable[1]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_data[33]~combout ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[14]~q ;
wire \jtag_uart_0|woverflow~q ;
wire \nios2_gen2_0|cpu|d_writedata[15]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~12_combout ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[15]~q ;
wire \jtag_uart_0|rvalid~q ;
wire \nios2_gen2_0|cpu|d_writedata[11]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~13_combout ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[11]~q ;
wire \nios2_gen2_0|cpu|d_writedata[13]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~14_combout ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[13]~q ;
wire \nios2_gen2_0|cpu|d_writedata[16]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~15_combout ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[16]~q ;
wire \jtag_uart_0|the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ;
wire \nios2_gen2_0|cpu|d_writedata[12]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~16_combout ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[12]~q ;
wire \jtag_uart_0|the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[27]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[28]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[29]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[30]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[31]~q ;
wire \nios2_gen2_0|cpu|d_writedata[10]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~17_combout ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[10]~q ;
wire \jtag_uart_0|ac~q ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[9]~q ;
wire \uart_0|the_processor_uart_0_regs|readdata[9]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~18_combout ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[8]~q ;
wire \uart_0|the_processor_uart_0_regs|readdata[8]~q ;
wire \nios2_gen2_0|cpu|d_writedata[8]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~19_combout ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[7]~q ;
wire \jtag_uart_0|av_readdata[7]~7_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~20_combout ;
wire \seg|readdata[7]~combout ;
wire \uart_0|the_processor_uart_0_regs|readdata[7]~q ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[6]~q ;
wire \jtag_uart_0|av_readdata[6]~8_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~21_combout ;
wire \seg|readdata[6]~combout ;
wire \uart_0|the_processor_uart_0_regs|readdata[6]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~2_combout ;
wire \nios2_gen2_0|cpu|d_writedata[21]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~22_combout ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[21]~q ;
wire \jtag_uart_0|the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ;
wire \nios2_gen2_0|cpu|d_writedata[20]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~23_combout ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[20]~q ;
wire \jtag_uart_0|the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~4_combout ;
wire \nios2_gen2_0|cpu|d_writedata[19]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~24_combout ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[19]~q ;
wire \jtag_uart_0|the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~6_combout ;
wire \nios2_gen2_0|cpu|d_writedata[18]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~25_combout ;
wire \jtag_uart_0|the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[18]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~8_combout ;
wire \nios2_gen2_0|cpu|d_writedata[17]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~26_combout ;
wire \jtag_uart_0|the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[17]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~10_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~11_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~13_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[9]~8_combout ;
wire \mm_interconnect_0|uart_0_s1_translator|end_begintransfer~q ;
wire \mm_interconnect_0|cmd_mux|src_data[38]~combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~0_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~0_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~1_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[38]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[39]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[40]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[41]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[42]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[43]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[44]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[45]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[32]~combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~1_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~2_combout ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[27]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~27_combout ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[28]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~28_combout ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[29]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~29_combout ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[30]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~30_combout ;
wire \nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[31]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~31_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~14_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~16_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~18_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~20_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~22_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~24_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~26_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~2_combout ;
wire \mm_interconnect_0|cmd_mux_007|src_payload~9_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~3_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~4_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~5_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[34]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~6_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~7_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[35]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~8_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~9_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~10_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~11_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~12_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[33]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~13_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~14_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~15_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~16_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~17_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~18_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~19_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~20_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~21_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~22_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~23_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~24_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~25_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~26_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~27_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~3_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~28_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~29_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~30_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~31_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~32_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~4_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~5_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~6_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~7_combout ;
wire \rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ;
wire \~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~8_combout ;
wire \auto_hub|~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ;
wire \clk_clk~input_o ;
wire \sw_export~input_o ;
wire \reset_reset_n~input_o ;
wire \uart_0_rxd~input_o ;
wire \altera_reserved_tms~input_o ;
wire \altera_reserved_tck~input_o ;
wire \altera_reserved_tdi~input_o ;
wire \altera_internal_jtag~TCKUTAP ;
wire \altera_internal_jtag~TMSUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ;
wire \altera_internal_jtag~TDIUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~16_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~15_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~15_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~16_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~6 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~8 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~10 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~12 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~12 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~23_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~17 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~19 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~15_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~22_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~19_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~15_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~17_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~18_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~16_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ;
wire \altera_internal_jtag~TDO ;


processor_processor_nios2_gen2_0 nios2_gen2_0(
	.sr_0(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[0]~q ),
	.W_alu_result_7(\nios2_gen2_0|cpu|W_alu_result[7]~q ),
	.W_alu_result_16(\nios2_gen2_0|cpu|W_alu_result[16]~q ),
	.W_alu_result_15(\nios2_gen2_0|cpu|W_alu_result[15]~q ),
	.W_alu_result_14(\nios2_gen2_0|cpu|W_alu_result[14]~q ),
	.W_alu_result_13(\nios2_gen2_0|cpu|W_alu_result[13]~q ),
	.W_alu_result_12(\nios2_gen2_0|cpu|W_alu_result[12]~q ),
	.W_alu_result_11(\nios2_gen2_0|cpu|W_alu_result[11]~q ),
	.W_alu_result_10(\nios2_gen2_0|cpu|W_alu_result[10]~q ),
	.W_alu_result_9(\nios2_gen2_0|cpu|W_alu_result[9]~q ),
	.W_alu_result_8(\nios2_gen2_0|cpu|W_alu_result[8]~q ),
	.W_alu_result_4(\nios2_gen2_0|cpu|W_alu_result[4]~q ),
	.W_alu_result_5(\nios2_gen2_0|cpu|W_alu_result[5]~q ),
	.W_alu_result_6(\nios2_gen2_0|cpu|W_alu_result[6]~q ),
	.W_alu_result_2(\nios2_gen2_0|cpu|W_alu_result[2]~q ),
	.W_alu_result_3(\nios2_gen2_0|cpu|W_alu_result[3]~q ),
	.q_a_22(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[22] ),
	.av_readdata_pre_22(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[22]~q ),
	.q_a_23(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_24(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[24] ),
	.q_a_25(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[25] ),
	.q_a_26(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[26] ),
	.q_a_1(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[1] ),
	.q_a_4(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[4] ),
	.q_a_3(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[3] ),
	.q_a_2(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[2] ),
	.q_a_5(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_14(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_15(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_13(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_16(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[16] ),
	.av_readdata_pre_16(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[16]~q ),
	.q_a_12(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_10(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_9(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_8(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_7(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[7] ),
	.q_a_6(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[6] ),
	.q_a_21(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[21] ),
	.av_readdata_pre_21(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[21]~q ),
	.q_a_20(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[20] ),
	.av_readdata_pre_20(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[20]~q ),
	.q_a_19(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[19] ),
	.av_readdata_pre_19(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[19]~q ),
	.q_a_18(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[18] ),
	.av_readdata_pre_18(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[18]~q ),
	.q_a_17(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[17] ),
	.av_readdata_pre_17(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[17]~q ),
	.readdata_0(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[0]~q ),
	.d_writedata_24(\nios2_gen2_0|cpu|d_writedata[24]~q ),
	.d_writedata_25(\nios2_gen2_0|cpu|d_writedata[25]~q ),
	.d_writedata_26(\nios2_gen2_0|cpu|d_writedata[26]~q ),
	.readdata_1(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[1]~q ),
	.readdata_3(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[3]~q ),
	.readdata_2(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[2]~q ),
	.q_a_27(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[27] ),
	.q_a_28(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[28] ),
	.q_a_29(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[29] ),
	.q_a_30(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[30] ),
	.q_a_31(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[31] ),
	.d_writedata_27(\nios2_gen2_0|cpu|d_writedata[27]~q ),
	.d_writedata_28(\nios2_gen2_0|cpu|d_writedata[28]~q ),
	.d_writedata_29(\nios2_gen2_0|cpu|d_writedata[29]~q ),
	.d_writedata_30(\nios2_gen2_0|cpu|d_writedata[30]~q ),
	.d_writedata_31(\nios2_gen2_0|cpu|d_writedata[31]~q ),
	.ir_out_0(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_tck|ir_out[0]~q ),
	.ir_out_1(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_tck|ir_out[1]~q ),
	.d_writedata_0(\nios2_gen2_0|cpu|d_writedata[0]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.d_write(\nios2_gen2_0|cpu|d_write~q ),
	.i_read(\nios2_gen2_0|cpu|i_read~q ),
	.F_pc_5(\nios2_gen2_0|cpu|F_pc[5]~q ),
	.F_pc_14(\nios2_gen2_0|cpu|F_pc[14]~q ),
	.F_pc_13(\nios2_gen2_0|cpu|F_pc[13]~q ),
	.F_pc_12(\nios2_gen2_0|cpu|F_pc[12]~q ),
	.F_pc_11(\nios2_gen2_0|cpu|F_pc[11]~q ),
	.F_pc_10(\nios2_gen2_0|cpu|F_pc[10]~q ),
	.F_pc_9(\nios2_gen2_0|cpu|F_pc[9]~q ),
	.F_pc_8(\nios2_gen2_0|cpu|F_pc[8]~q ),
	.F_pc_7(\nios2_gen2_0|cpu|F_pc[7]~q ),
	.F_pc_6(\nios2_gen2_0|cpu|F_pc[6]~q ),
	.F_pc_2(\nios2_gen2_0|cpu|F_pc[2]~q ),
	.F_pc_3(\nios2_gen2_0|cpu|F_pc[3]~q ),
	.F_pc_4(\nios2_gen2_0|cpu|F_pc[4]~q ),
	.d_read(\nios2_gen2_0|cpu|d_read~q ),
	.F_pc_1(\nios2_gen2_0|cpu|F_pc[1]~q ),
	.F_pc_0(\nios2_gen2_0|cpu|F_pc[0]~q ),
	.d_writedata_1(\nios2_gen2_0|cpu|d_writedata[1]~q ),
	.d_writedata_2(\nios2_gen2_0|cpu|d_writedata[2]~q ),
	.d_writedata_3(\nios2_gen2_0|cpu|d_writedata[3]~q ),
	.d_writedata_4(\nios2_gen2_0|cpu|d_writedata[4]~q ),
	.d_writedata_5(\nios2_gen2_0|cpu|d_writedata[5]~q ),
	.d_writedata_6(\nios2_gen2_0|cpu|d_writedata[6]~q ),
	.d_writedata_7(\nios2_gen2_0|cpu|d_writedata[7]~q ),
	.src0_valid(\mm_interconnect_0|rsp_demux|src0_valid~0_combout ),
	.read_latency_shift_reg_0(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|mem[0][56]~q ),
	.src0_valid1(\mm_interconnect_0|rsp_demux_001|src0_valid~0_combout ),
	.read_latency_shift_reg_01(\mm_interconnect_0|onchip_memory2_0_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_74_01(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_01(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][56]~q ),
	.src0_valid2(\mm_interconnect_0|rsp_demux_002|src0_valid~0_combout ),
	.src0_valid3(\mm_interconnect_0|rsp_demux_003|src0_valid~0_combout ),
	.WideOr1(\mm_interconnect_0|rsp_mux|WideOr1~0_combout ),
	.src0_valid4(\mm_interconnect_0|rsp_demux_004|src0_valid~0_combout ),
	.read_latency_shift_reg_02(\mm_interconnect_0|seg_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_74_02(\mm_interconnect_0|seg_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_02(\mm_interconnect_0|seg_s1_agent_rsp_fifo|mem[0][56]~q ),
	.src0_valid5(\mm_interconnect_0|rsp_demux_005|src0_valid~0_combout ),
	.src0_valid6(\mm_interconnect_0|rsp_demux_007|src0_valid~0_combout ),
	.WideOr11(\mm_interconnect_0|rsp_mux|WideOr1~1_combout ),
	.WideOr12(\mm_interconnect_0|rsp_mux|WideOr1~combout ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_001|saved_grant[0]~q ),
	.debug_mem_slave_waitrequest(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|the_processor_nios2_gen2_0_cpu_nios2_ocimem|waitrequest~q ),
	.mem_used_1(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|mem_used[1]~q ),
	.av_waitrequest(\mm_interconnect_0|nios2_gen2_0_data_master_translator|av_waitrequest~1_combout ),
	.src1_valid(\mm_interconnect_0|rsp_demux|src1_valid~0_combout ),
	.src1_valid1(\mm_interconnect_0|rsp_demux_001|src1_valid~0_combout ),
	.src1_valid2(\mm_interconnect_0|rsp_demux_002|src1_valid~0_combout ),
	.src1_valid3(\mm_interconnect_0|rsp_demux_005|src1_valid~0_combout ),
	.WideOr13(\mm_interconnect_0|rsp_mux_001|WideOr1~0_combout ),
	.src1_valid4(\mm_interconnect_0|rsp_demux_007|src1_valid~0_combout ),
	.src_payload(\mm_interconnect_0|rsp_mux_001|src_payload~0_combout ),
	.src_payload1(\mm_interconnect_0|rsp_mux_001|src_payload~1_combout ),
	.WideOr14(\mm_interconnect_0|rsp_mux_001|WideOr1~1_combout ),
	.uav_write(\mm_interconnect_0|nios2_gen2_0_data_master_translator|uav_write~0_combout ),
	.d_writedata_9(\nios2_gen2_0|cpu|d_writedata[9]~q ),
	.WideOr15(\mm_interconnect_0|cmd_mux_001|WideOr1~combout ),
	.rf_source_valid(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_agent|rf_source_valid~0_combout ),
	.hbreak_enabled(\nios2_gen2_0|cpu|hbreak_enabled~q ),
	.src_data_0(\mm_interconnect_0|rsp_mux|src_data[0]~combout ),
	.av_readdata_pre_221(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[22]~q ),
	.av_readdata_pre_23(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[23]~q ),
	.av_readdata_pre_24(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[24]~q ),
	.av_readdata_pre_25(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[25]~q ),
	.av_readdata_pre_26(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[26]~q ),
	.src_data_01(\mm_interconnect_0|rsp_mux_001|src_data[0]~0_combout ),
	.src_data_02(\mm_interconnect_0|rsp_mux_001|src_data[0]~1_combout ),
	.src_data_03(\mm_interconnect_0|rsp_mux_001|src_data[0]~3_combout ),
	.av_readdata_pre_1(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_11(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_12(\mm_interconnect_0|uart_0_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_13(\mm_interconnect_0|seg_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_14(\mm_interconnect_0|led_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_15(\mm_interconnect_0|seg_en_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_4(\mm_interconnect_0|seg_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_41(\mm_interconnect_0|uart_0_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_42(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_43(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_3(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[3]~q ),
	.src_payload2(\mm_interconnect_0|rsp_mux_001|src_payload~4_combout ),
	.av_readdata_pre_31(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_32(\mm_interconnect_0|uart_0_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_33(\mm_interconnect_0|seg_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_2(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_27(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_28(\mm_interconnect_0|seg_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_29(\mm_interconnect_0|seg_en_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_210(\mm_interconnect_0|uart_0_s1_translator|av_readdata_pre[2]~q ),
	.src_data_46(\mm_interconnect_0|cmd_mux_001|src_data[46]~combout ),
	.av_readdata_pre_5(\mm_interconnect_0|seg_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_51(\mm_interconnect_0|uart_0_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_52(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_53(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_141(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_142(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_151(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_152(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[15]~q ),
	.src_payload3(\mm_interconnect_0|rsp_mux_001|src_payload~5_combout ),
	.av_readdata_pre_111(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[11]~q ),
	.av_readdata_pre_131(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_132(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_161(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[16]~q ),
	.av_readdata_pre_121(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_122(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_10(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_101(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_9(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_91(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_92(\mm_interconnect_0|uart_0_s1_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_8(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_81(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_82(\mm_interconnect_0|uart_0_s1_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_7(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_71(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_72(\mm_interconnect_0|seg_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_73(\mm_interconnect_0|uart_0_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_6(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_61(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_62(\mm_interconnect_0|seg_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_63(\mm_interconnect_0|uart_0_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_211(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_201(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_191(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[19]~q ),
	.av_readdata_pre_181(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_171(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[17]~q ),
	.r_early_rst(\rst_controller|r_early_rst~q ),
	.src_data_8(\mm_interconnect_0|rsp_mux|src_data[8]~5_combout ),
	.d_byteenable_0(\nios2_gen2_0|cpu|d_byteenable[0]~q ),
	.av_readdata_9(\jtag_uart_0|av_readdata[9]~combout ),
	.av_readdata_8(\jtag_uart_0|av_readdata[8]~1_combout ),
	.irq(\uart_0|the_processor_uart_0_regs|irq~q ),
	.d_writedata_22(\nios2_gen2_0|cpu|d_writedata[22]~q ),
	.d_byteenable_2(\nios2_gen2_0|cpu|d_byteenable[2]~q ),
	.readdata_22(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[22]~q ),
	.readdata_23(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[23]~q ),
	.d_writedata_23(\nios2_gen2_0|cpu|d_writedata[23]~q ),
	.readdata_24(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[24]~q ),
	.d_byteenable_3(\nios2_gen2_0|cpu|d_byteenable[3]~q ),
	.readdata_25(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[25]~q ),
	.readdata_26(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[26]~q ),
	.readdata_4(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[4]~q ),
	.readdata_5(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[5]~q ),
	.d_writedata_14(\nios2_gen2_0|cpu|d_writedata[14]~q ),
	.d_byteenable_1(\nios2_gen2_0|cpu|d_byteenable[1]~q ),
	.readdata_14(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[14]~q ),
	.d_writedata_15(\nios2_gen2_0|cpu|d_writedata[15]~q ),
	.readdata_15(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[15]~q ),
	.d_writedata_11(\nios2_gen2_0|cpu|d_writedata[11]~q ),
	.readdata_11(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[11]~q ),
	.d_writedata_13(\nios2_gen2_0|cpu|d_writedata[13]~q ),
	.readdata_13(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[13]~q ),
	.d_writedata_16(\nios2_gen2_0|cpu|d_writedata[16]~q ),
	.readdata_16(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[16]~q ),
	.d_writedata_12(\nios2_gen2_0|cpu|d_writedata[12]~q ),
	.readdata_12(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[12]~q ),
	.av_readdata_pre_271(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[27]~q ),
	.av_readdata_pre_281(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[28]~q ),
	.av_readdata_pre_291(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[29]~q ),
	.av_readdata_pre_30(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[30]~q ),
	.av_readdata_pre_311(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[31]~q ),
	.d_writedata_10(\nios2_gen2_0|cpu|d_writedata[10]~q ),
	.readdata_10(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[10]~q ),
	.readdata_9(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[9]~q ),
	.readdata_8(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[8]~q ),
	.d_writedata_8(\nios2_gen2_0|cpu|d_writedata[8]~q ),
	.readdata_7(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[7]~q ),
	.readdata_6(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[6]~q ),
	.src_payload4(\mm_interconnect_0|rsp_mux|src_payload~2_combout ),
	.d_writedata_21(\nios2_gen2_0|cpu|d_writedata[21]~q ),
	.readdata_21(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[21]~q ),
	.d_writedata_20(\nios2_gen2_0|cpu|d_writedata[20]~q ),
	.readdata_20(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[20]~q ),
	.src_payload5(\mm_interconnect_0|rsp_mux|src_payload~4_combout ),
	.d_writedata_19(\nios2_gen2_0|cpu|d_writedata[19]~q ),
	.readdata_19(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[19]~q ),
	.src_payload6(\mm_interconnect_0|rsp_mux|src_payload~6_combout ),
	.d_writedata_18(\nios2_gen2_0|cpu|d_writedata[18]~q ),
	.readdata_18(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[18]~q ),
	.src_payload7(\mm_interconnect_0|rsp_mux|src_payload~8_combout ),
	.d_writedata_17(\nios2_gen2_0|cpu|d_writedata[17]~q ),
	.readdata_17(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[17]~q ),
	.src_payload8(\mm_interconnect_0|rsp_mux|src_payload~10_combout ),
	.src_payload9(\mm_interconnect_0|rsp_mux|src_payload~11_combout ),
	.src_payload10(\mm_interconnect_0|rsp_mux|src_payload~13_combout ),
	.src_data_9(\mm_interconnect_0|rsp_mux|src_data[9]~8_combout ),
	.src_payload11(\mm_interconnect_0|cmd_mux_001|src_payload~0_combout ),
	.src_payload12(\mm_interconnect_0|cmd_mux_001|src_payload~1_combout ),
	.src_data_38(\mm_interconnect_0|cmd_mux_001|src_data[38]~combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux_001|src_data[39]~combout ),
	.src_data_40(\mm_interconnect_0|cmd_mux_001|src_data[40]~combout ),
	.src_data_41(\mm_interconnect_0|cmd_mux_001|src_data[41]~combout ),
	.src_data_42(\mm_interconnect_0|cmd_mux_001|src_data[42]~combout ),
	.src_data_43(\mm_interconnect_0|cmd_mux_001|src_data[43]~combout ),
	.src_data_44(\mm_interconnect_0|cmd_mux_001|src_data[44]~combout ),
	.src_data_45(\mm_interconnect_0|cmd_mux_001|src_data[45]~combout ),
	.src_data_32(\mm_interconnect_0|cmd_mux_001|src_data[32]~combout ),
	.readdata_27(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[27]~q ),
	.readdata_28(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[28]~q ),
	.readdata_29(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[29]~q ),
	.readdata_30(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[30]~q ),
	.readdata_31(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[31]~q ),
	.src_payload13(\mm_interconnect_0|rsp_mux|src_payload~14_combout ),
	.src_payload14(\mm_interconnect_0|rsp_mux|src_payload~16_combout ),
	.src_payload15(\mm_interconnect_0|rsp_mux|src_payload~18_combout ),
	.src_payload16(\mm_interconnect_0|rsp_mux|src_payload~20_combout ),
	.src_payload17(\mm_interconnect_0|rsp_mux|src_payload~22_combout ),
	.src_payload18(\mm_interconnect_0|rsp_mux|src_payload~24_combout ),
	.src_payload19(\mm_interconnect_0|rsp_mux|src_payload~26_combout ),
	.src_payload20(\mm_interconnect_0|cmd_mux_001|src_payload~2_combout ),
	.src_payload21(\mm_interconnect_0|cmd_mux_001|src_payload~3_combout ),
	.src_payload22(\mm_interconnect_0|cmd_mux_001|src_payload~4_combout ),
	.src_payload23(\mm_interconnect_0|cmd_mux_001|src_payload~5_combout ),
	.src_data_34(\mm_interconnect_0|cmd_mux_001|src_data[34]~combout ),
	.src_payload24(\mm_interconnect_0|cmd_mux_001|src_payload~6_combout ),
	.src_payload25(\mm_interconnect_0|cmd_mux_001|src_payload~7_combout ),
	.src_data_35(\mm_interconnect_0|cmd_mux_001|src_data[35]~combout ),
	.src_payload26(\mm_interconnect_0|cmd_mux_001|src_payload~8_combout ),
	.src_payload27(\mm_interconnect_0|cmd_mux_001|src_payload~9_combout ),
	.src_payload28(\mm_interconnect_0|cmd_mux_001|src_payload~10_combout ),
	.src_payload29(\mm_interconnect_0|cmd_mux_001|src_payload~11_combout ),
	.src_payload30(\mm_interconnect_0|cmd_mux_001|src_payload~12_combout ),
	.src_data_33(\mm_interconnect_0|cmd_mux_001|src_data[33]~combout ),
	.src_payload31(\mm_interconnect_0|cmd_mux_001|src_payload~13_combout ),
	.src_payload32(\mm_interconnect_0|cmd_mux_001|src_payload~14_combout ),
	.src_payload33(\mm_interconnect_0|cmd_mux_001|src_payload~15_combout ),
	.src_payload34(\mm_interconnect_0|cmd_mux_001|src_payload~16_combout ),
	.src_payload35(\mm_interconnect_0|cmd_mux_001|src_payload~17_combout ),
	.src_payload36(\mm_interconnect_0|cmd_mux_001|src_payload~18_combout ),
	.src_payload37(\mm_interconnect_0|cmd_mux_001|src_payload~19_combout ),
	.src_payload38(\mm_interconnect_0|cmd_mux_001|src_payload~20_combout ),
	.src_payload39(\mm_interconnect_0|cmd_mux_001|src_payload~21_combout ),
	.src_payload40(\mm_interconnect_0|cmd_mux_001|src_payload~22_combout ),
	.src_payload41(\mm_interconnect_0|cmd_mux_001|src_payload~23_combout ),
	.src_payload42(\mm_interconnect_0|cmd_mux_001|src_payload~24_combout ),
	.src_payload43(\mm_interconnect_0|cmd_mux_001|src_payload~25_combout ),
	.src_payload44(\mm_interconnect_0|cmd_mux_001|src_payload~26_combout ),
	.src_payload45(\mm_interconnect_0|cmd_mux_001|src_payload~27_combout ),
	.src_payload46(\mm_interconnect_0|cmd_mux_001|src_payload~28_combout ),
	.src_payload47(\mm_interconnect_0|cmd_mux_001|src_payload~29_combout ),
	.src_payload48(\mm_interconnect_0|cmd_mux_001|src_payload~30_combout ),
	.src_payload49(\mm_interconnect_0|cmd_mux_001|src_payload~31_combout ),
	.src_payload50(\mm_interconnect_0|cmd_mux_001|src_payload~32_combout ),
	.altera_internal_jtag(\altera_internal_jtag~TCKUTAP ),
	.altera_internal_jtag1(\altera_internal_jtag~TDIUTAP ),
	.state_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.state_4(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.virtual_ir_scan_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.state_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.state_8(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.splitter_nodes_receive_1_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ),
	.irf_reg_0_2(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.irf_reg_1_2(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.clk_clk(\clk_clk~input_o ));

processor_processor_mm_interconnect_0 mm_interconnect_0(
	.W_alu_result_7(\nios2_gen2_0|cpu|W_alu_result[7]~q ),
	.W_alu_result_16(\nios2_gen2_0|cpu|W_alu_result[16]~q ),
	.W_alu_result_15(\nios2_gen2_0|cpu|W_alu_result[15]~q ),
	.W_alu_result_14(\nios2_gen2_0|cpu|W_alu_result[14]~q ),
	.W_alu_result_13(\nios2_gen2_0|cpu|W_alu_result[13]~q ),
	.W_alu_result_12(\nios2_gen2_0|cpu|W_alu_result[12]~q ),
	.W_alu_result_11(\nios2_gen2_0|cpu|W_alu_result[11]~q ),
	.W_alu_result_10(\nios2_gen2_0|cpu|W_alu_result[10]~q ),
	.W_alu_result_9(\nios2_gen2_0|cpu|W_alu_result[9]~q ),
	.W_alu_result_8(\nios2_gen2_0|cpu|W_alu_result[8]~q ),
	.W_alu_result_4(\nios2_gen2_0|cpu|W_alu_result[4]~q ),
	.W_alu_result_5(\nios2_gen2_0|cpu|W_alu_result[5]~q ),
	.W_alu_result_6(\nios2_gen2_0|cpu|W_alu_result[6]~q ),
	.W_alu_result_2(\nios2_gen2_0|cpu|W_alu_result[2]~q ),
	.W_alu_result_3(\nios2_gen2_0|cpu|W_alu_result[3]~q ),
	.q_a_0(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[0] ),
	.q_a_22(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[22] ),
	.av_readdata_pre_22(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[22]~q ),
	.q_a_23(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_14(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_15(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_11(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_13(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_16(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[16] ),
	.av_readdata_pre_16(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[16]~q ),
	.q_a_12(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_10(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_9(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_8(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_21(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[21] ),
	.av_readdata_pre_21(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[21]~q ),
	.q_a_20(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[20] ),
	.av_readdata_pre_20(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[20]~q ),
	.q_a_19(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[19] ),
	.av_readdata_pre_19(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[19]~q ),
	.q_a_18(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[18] ),
	.av_readdata_pre_18(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[18]~q ),
	.q_a_17(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[17] ),
	.av_readdata_pre_17(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[17]~q ),
	.readdata_0(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[0]~q ),
	.d_writedata_24(\nios2_gen2_0|cpu|d_writedata[24]~q ),
	.d_writedata_25(\nios2_gen2_0|cpu|d_writedata[25]~q ),
	.d_writedata_26(\nios2_gen2_0|cpu|d_writedata[26]~q ),
	.readdata_1(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[1]~q ),
	.readdata_3(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[3]~q ),
	.readdata_2(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[2]~q ),
	.d_writedata_27(\nios2_gen2_0|cpu|d_writedata[27]~q ),
	.d_writedata_28(\nios2_gen2_0|cpu|d_writedata[28]~q ),
	.d_writedata_29(\nios2_gen2_0|cpu|d_writedata[29]~q ),
	.d_writedata_30(\nios2_gen2_0|cpu|d_writedata[30]~q ),
	.d_writedata_31(\nios2_gen2_0|cpu|d_writedata[31]~q ),
	.d_writedata_0(\nios2_gen2_0|cpu|d_writedata[0]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_003|saved_grant[0]~q ),
	.d_write(\nios2_gen2_0|cpu|d_write~q ),
	.src_payload(\mm_interconnect_0|cmd_mux_003|src_payload~0_combout ),
	.saved_grant_1(\mm_interconnect_0|cmd_mux_003|saved_grant[1]~q ),
	.rst1(\jtag_uart_0|processor_jtag_uart_0_alt_jtag_atlantic|rst1~q ),
	.i_read(\nios2_gen2_0|cpu|i_read~q ),
	.F_pc_5(\nios2_gen2_0|cpu|F_pc[5]~q ),
	.F_pc_14(\nios2_gen2_0|cpu|F_pc[14]~q ),
	.F_pc_13(\nios2_gen2_0|cpu|F_pc[13]~q ),
	.F_pc_12(\nios2_gen2_0|cpu|F_pc[12]~q ),
	.F_pc_11(\nios2_gen2_0|cpu|F_pc[11]~q ),
	.F_pc_10(\nios2_gen2_0|cpu|F_pc[10]~q ),
	.F_pc_9(\nios2_gen2_0|cpu|F_pc[9]~q ),
	.F_pc_8(\nios2_gen2_0|cpu|F_pc[8]~q ),
	.F_pc_7(\nios2_gen2_0|cpu|F_pc[7]~q ),
	.F_pc_6(\nios2_gen2_0|cpu|F_pc[6]~q ),
	.F_pc_2(\nios2_gen2_0|cpu|F_pc[2]~q ),
	.F_pc_3(\nios2_gen2_0|cpu|F_pc[3]~q ),
	.F_pc_4(\nios2_gen2_0|cpu|F_pc[4]~q ),
	.src_valid(\mm_interconnect_0|cmd_mux_003|src_valid~3_combout ),
	.d_read(\nios2_gen2_0|cpu|d_read~q ),
	.src_valid1(\mm_interconnect_0|cmd_mux_003|src_valid~5_combout ),
	.mem_used_1(\mm_interconnect_0|led_s1_agent_rsp_fifo|mem_used[1]~q ),
	.always0(\led|always0~0_combout ),
	.F_pc_1(\nios2_gen2_0|cpu|F_pc[1]~q ),
	.F_pc_0(\nios2_gen2_0|cpu|F_pc[0]~q ),
	.wait_latency_counter_1(\mm_interconnect_0|led_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|led_s1_translator|wait_latency_counter[0]~q ),
	.d_writedata_1(\nios2_gen2_0|cpu|d_writedata[1]~q ),
	.saved_grant_01(\mm_interconnect_0|cmd_mux_005|saved_grant[0]~q ),
	.src_payload1(\mm_interconnect_0|cmd_mux_005|src_payload~0_combout ),
	.saved_grant_11(\mm_interconnect_0|cmd_mux_005|saved_grant[1]~q ),
	.src_valid2(\mm_interconnect_0|cmd_mux_005|src_valid~2_combout ),
	.src_valid3(\mm_interconnect_0|cmd_mux_005|src_valid~4_combout ),
	.mem_used_11(\mm_interconnect_0|seg_s1_agent_rsp_fifo|mem_used[1]~q ),
	.always01(\seg|always0~0_combout ),
	.wait_latency_counter_11(\mm_interconnect_0|seg_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_01(\mm_interconnect_0|seg_s1_translator|wait_latency_counter[0]~q ),
	.d_writedata_2(\nios2_gen2_0|cpu|d_writedata[2]~q ),
	.d_writedata_3(\nios2_gen2_0|cpu|d_writedata[3]~q ),
	.d_writedata_4(\nios2_gen2_0|cpu|d_writedata[4]~q ),
	.d_writedata_5(\nios2_gen2_0|cpu|d_writedata[5]~q ),
	.d_writedata_6(\nios2_gen2_0|cpu|d_writedata[6]~q ),
	.d_writedata_7(\nios2_gen2_0|cpu|d_writedata[7]~q ),
	.saved_grant_02(\mm_interconnect_0|cmd_mux_004|saved_grant[0]~q ),
	.src_payload2(\mm_interconnect_0|cmd_mux_004|src_payload~0_combout ),
	.saved_grant_12(\mm_interconnect_0|cmd_mux_004|saved_grant[1]~q ),
	.src_valid4(\mm_interconnect_0|cmd_mux_004|src_valid~3_combout ),
	.src_valid5(\mm_interconnect_0|cmd_mux_004|src_valid~5_combout ),
	.mem_used_12(\mm_interconnect_0|seg_en_s1_agent_rsp_fifo|mem_used[1]~q ),
	.always02(\seg_en|always0~0_combout ),
	.wait_latency_counter_12(\mm_interconnect_0|seg_en_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_02(\mm_interconnect_0|seg_en_s1_translator|wait_latency_counter[0]~q ),
	.src0_valid(\mm_interconnect_0|rsp_demux|src0_valid~0_combout ),
	.read_latency_shift_reg_0(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|mem[0][56]~q ),
	.src0_valid1(\mm_interconnect_0|rsp_demux_001|src0_valid~0_combout ),
	.read_latency_shift_reg_01(\mm_interconnect_0|onchip_memory2_0_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_74_01(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_01(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][56]~q ),
	.src0_valid2(\mm_interconnect_0|rsp_demux_002|src0_valid~0_combout ),
	.src0_valid3(\mm_interconnect_0|rsp_demux_003|src0_valid~0_combout ),
	.WideOr1(\mm_interconnect_0|rsp_mux|WideOr1~0_combout ),
	.src0_valid4(\mm_interconnect_0|rsp_demux_004|src0_valid~0_combout ),
	.read_latency_shift_reg_02(\mm_interconnect_0|seg_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_74_02(\mm_interconnect_0|seg_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_02(\mm_interconnect_0|seg_s1_agent_rsp_fifo|mem[0][56]~q ),
	.src0_valid5(\mm_interconnect_0|rsp_demux_005|src0_valid~0_combout ),
	.src0_valid6(\mm_interconnect_0|rsp_demux_007|src0_valid~0_combout ),
	.WideOr11(\mm_interconnect_0|rsp_mux|WideOr1~1_combout ),
	.WideOr12(\mm_interconnect_0|rsp_mux|WideOr1~combout ),
	.saved_grant_03(\mm_interconnect_0|cmd_mux_002|saved_grant[0]~q ),
	.mem_used_13(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem_used[1]~q ),
	.mem_used_14(\mm_interconnect_0|uart_0_s1_agent_rsp_fifo|mem_used[1]~q ),
	.wait_latency_counter_13(\mm_interconnect_0|uart_0_s1_translator|wait_latency_counter[1]~q ),
	.av_waitrequest(\jtag_uart_0|av_waitrequest~q ),
	.mem_used_15(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo|mem_used[1]~q ),
	.saved_grant_04(\mm_interconnect_0|cmd_mux|saved_grant[0]~q ),
	.saved_grant_05(\mm_interconnect_0|cmd_mux_001|saved_grant[0]~q ),
	.waitrequest(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|the_processor_nios2_gen2_0_cpu_nios2_ocimem|waitrequest~q ),
	.mem_used_16(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|mem_used[1]~q ),
	.saved_grant_06(\mm_interconnect_0|cmd_mux_006|saved_grant[0]~q ),
	.saved_grant_13(\mm_interconnect_0|cmd_mux_006|saved_grant[1]~q ),
	.nios2_gen2_0_data_master_waitrequest(\mm_interconnect_0|nios2_gen2_0_data_master_translator|av_waitrequest~1_combout ),
	.src1_valid(\mm_interconnect_0|rsp_demux|src1_valid~0_combout ),
	.src1_valid1(\mm_interconnect_0|rsp_demux_001|src1_valid~0_combout ),
	.src1_valid2(\mm_interconnect_0|rsp_demux_002|src1_valid~0_combout ),
	.src1_valid3(\mm_interconnect_0|rsp_demux_005|src1_valid~0_combout ),
	.WideOr13(\mm_interconnect_0|rsp_mux_001|WideOr1~0_combout ),
	.src1_valid4(\mm_interconnect_0|rsp_demux_007|src1_valid~0_combout ),
	.src_payload3(\mm_interconnect_0|rsp_mux_001|src_payload~0_combout ),
	.src_payload4(\mm_interconnect_0|rsp_mux_001|src_payload~1_combout ),
	.WideOr14(\mm_interconnect_0|rsp_mux_001|WideOr1~1_combout ),
	.uav_write(\mm_interconnect_0|nios2_gen2_0_data_master_translator|uav_write~0_combout ),
	.d_writedata_9(\nios2_gen2_0|cpu|d_writedata[9]~q ),
	.src_payload5(\mm_interconnect_0|cmd_mux_007|src_payload~0_combout ),
	.src_data_38(\mm_interconnect_0|cmd_mux_007|src_data[38]~combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux_007|src_data[39]~combout ),
	.src_data_40(\mm_interconnect_0|cmd_mux_007|src_data[40]~combout ),
	.WideOr15(\mm_interconnect_0|cmd_mux_007|WideOr1~combout ),
	.uart_0_s1_begintransfer(\mm_interconnect_0|uart_0_s1_translator|av_begintransfer~0_combout ),
	.src_data_56(\mm_interconnect_0|cmd_mux|src_data[56]~combout ),
	.WideOr16(\mm_interconnect_0|cmd_mux|WideOr1~combout ),
	.WideOr17(\mm_interconnect_0|cmd_mux_001|WideOr1~combout ),
	.WideOr18(\mm_interconnect_0|cmd_mux_002|WideOr1~combout ),
	.src_data_561(\mm_interconnect_0|cmd_mux_007|src_data[56]~combout ),
	.rx_rd_strobe_onset(\uart_0|the_processor_uart_0_rx|rx_rd_strobe_onset~0_combout ),
	.rf_source_valid(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_agent|rf_source_valid~0_combout ),
	.hbreak_enabled(\nios2_gen2_0|cpu|hbreak_enabled~q ),
	.src_data_0(\mm_interconnect_0|rsp_mux|src_data[0]~combout ),
	.av_readdata_pre_221(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[22]~q ),
	.av_readdata_pre_23(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[23]~q ),
	.av_readdata_pre_24(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[24]~q ),
	.av_readdata_pre_25(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[25]~q ),
	.av_readdata_pre_26(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[26]~q ),
	.src_data_01(\mm_interconnect_0|rsp_mux_001|src_data[0]~0_combout ),
	.src_data_02(\mm_interconnect_0|rsp_mux_001|src_data[0]~1_combout ),
	.src_data_03(\mm_interconnect_0|rsp_mux_001|src_data[0]~3_combout ),
	.av_readdata_pre_1(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_11(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_12(\mm_interconnect_0|uart_0_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_13(\mm_interconnect_0|seg_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_14(\mm_interconnect_0|led_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_15(\mm_interconnect_0|seg_en_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_4(\mm_interconnect_0|seg_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_41(\mm_interconnect_0|uart_0_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_42(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_43(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_3(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[3]~q ),
	.src_payload6(\mm_interconnect_0|rsp_mux_001|src_payload~4_combout ),
	.av_readdata_pre_31(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_32(\mm_interconnect_0|uart_0_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_33(\mm_interconnect_0|seg_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_2(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_27(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_28(\mm_interconnect_0|seg_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_29(\mm_interconnect_0|seg_en_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_210(\mm_interconnect_0|uart_0_s1_translator|av_readdata_pre[2]~q ),
	.src_data_46(\mm_interconnect_0|cmd_mux_001|src_data[46]~combout ),
	.av_readdata_pre_5(\mm_interconnect_0|seg_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_51(\mm_interconnect_0|uart_0_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_52(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_53(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_141(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_142(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_151(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_152(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[15]~q ),
	.src_payload7(\mm_interconnect_0|rsp_mux_001|src_payload~5_combout ),
	.av_readdata_pre_111(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[11]~q ),
	.av_readdata_pre_131(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_132(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_161(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[16]~q ),
	.av_readdata_pre_121(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_122(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_10(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_101(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_9(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_91(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_92(\mm_interconnect_0|uart_0_s1_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_8(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_81(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_82(\mm_interconnect_0|uart_0_s1_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_7(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_71(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_72(\mm_interconnect_0|seg_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_73(\mm_interconnect_0|uart_0_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_6(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_61(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_62(\mm_interconnect_0|seg_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_63(\mm_interconnect_0|uart_0_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_211(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_201(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_191(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[19]~q ),
	.av_readdata_pre_181(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_171(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[17]~q ),
	.src_payload8(\mm_interconnect_0|cmd_mux_007|src_payload~1_combout ),
	.src_payload9(\mm_interconnect_0|cmd_mux_007|src_payload~2_combout ),
	.src_payload10(\mm_interconnect_0|cmd_mux_007|src_payload~3_combout ),
	.src_payload11(\mm_interconnect_0|cmd_mux_007|src_payload~4_combout ),
	.src_payload12(\mm_interconnect_0|cmd_mux_007|src_payload~5_combout ),
	.src_payload13(\mm_interconnect_0|cmd_mux_007|src_payload~6_combout ),
	.src_payload14(\mm_interconnect_0|cmd_mux_007|src_payload~7_combout ),
	.src_payload15(\mm_interconnect_0|cmd_mux_007|src_payload~8_combout ),
	.b_full(\jtag_uart_0|the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.src_data_8(\mm_interconnect_0|rsp_mux|src_data[8]~5_combout ),
	.readdata_01(\seg|readdata[0]~combout ),
	.readdata_02(\seg_en|readdata[0]~combout ),
	.src_payload16(\mm_interconnect_0|cmd_mux_002|src_payload~0_combout ),
	.src_data_381(\mm_interconnect_0|cmd_mux_002|src_data[38]~combout ),
	.src_data_391(\mm_interconnect_0|cmd_mux_002|src_data[39]~combout ),
	.src_data_401(\mm_interconnect_0|cmd_mux_002|src_data[40]~combout ),
	.src_data_41(\mm_interconnect_0|cmd_mux_002|src_data[41]~combout ),
	.src_data_42(\mm_interconnect_0|cmd_mux_002|src_data[42]~combout ),
	.src_data_43(\mm_interconnect_0|cmd_mux_002|src_data[43]~combout ),
	.src_data_44(\mm_interconnect_0|cmd_mux_002|src_data[44]~combout ),
	.src_data_45(\mm_interconnect_0|cmd_mux_002|src_data[45]~combout ),
	.src_data_461(\mm_interconnect_0|cmd_mux_002|src_data[46]~combout ),
	.src_data_47(\mm_interconnect_0|cmd_mux_002|src_data[47]~combout ),
	.src_data_48(\mm_interconnect_0|cmd_mux_002|src_data[48]~combout ),
	.src_data_49(\mm_interconnect_0|cmd_mux_002|src_data[49]~combout ),
	.src_data_50(\mm_interconnect_0|cmd_mux_002|src_data[50]~combout ),
	.d_byteenable_0(\nios2_gen2_0|cpu|d_byteenable[0]~q ),
	.src_data_32(\mm_interconnect_0|cmd_mux_002|src_data[32]~combout ),
	.read_0(\jtag_uart_0|read_0~q ),
	.av_readdata_0(\jtag_uart_0|av_readdata[0]~0_combout ),
	.readdata_03(\uart_0|the_processor_uart_0_regs|readdata[0]~q ),
	.readdata_04(\led|readdata[0]~combout ),
	.readdata_05(\sw|readdata[0]~q ),
	.av_readdata_9(\jtag_uart_0|av_readdata[9]~combout ),
	.av_readdata_8(\jtag_uart_0|av_readdata[8]~1_combout ),
	.d_writedata_22(\nios2_gen2_0|cpu|d_writedata[22]~q ),
	.src_payload17(\mm_interconnect_0|cmd_mux_002|src_payload~1_combout ),
	.d_byteenable_2(\nios2_gen2_0|cpu|d_byteenable[2]~q ),
	.src_data_34(\mm_interconnect_0|cmd_mux_002|src_data[34]~combout ),
	.readdata_22(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[22]~q ),
	.b_full1(\jtag_uart_0|the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.counter_reg_bit_5(\jtag_uart_0|the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.counter_reg_bit_4(\jtag_uart_0|the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\jtag_uart_0|the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\jtag_uart_0|the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\jtag_uart_0|the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\jtag_uart_0|the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.readdata_23(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[23]~q ),
	.d_writedata_23(\nios2_gen2_0|cpu|d_writedata[23]~q ),
	.src_payload18(\mm_interconnect_0|cmd_mux_002|src_payload~2_combout ),
	.readdata_24(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[24]~q ),
	.src_payload19(\mm_interconnect_0|cmd_mux_002|src_payload~3_combout ),
	.d_byteenable_3(\nios2_gen2_0|cpu|d_byteenable[3]~q ),
	.src_data_35(\mm_interconnect_0|cmd_mux_002|src_data[35]~combout ),
	.readdata_25(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[25]~q ),
	.src_payload20(\mm_interconnect_0|cmd_mux_002|src_payload~4_combout ),
	.readdata_26(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[26]~q ),
	.src_payload21(\mm_interconnect_0|cmd_mux_002|src_payload~5_combout ),
	.av_readdata_1(\jtag_uart_0|av_readdata[1]~2_combout ),
	.src_payload22(\mm_interconnect_0|cmd_mux_002|src_payload~6_combout ),
	.readdata_11(\uart_0|the_processor_uart_0_regs|readdata[1]~q ),
	.readdata_12(\seg|readdata[1]~combout ),
	.readdata_13(\led|readdata[1]~combout ),
	.readdata_14(\seg_en|readdata[1]~combout ),
	.src_payload23(\mm_interconnect_0|cmd_mux_002|src_payload~7_combout ),
	.readdata_4(\seg|readdata[4]~combout ),
	.readdata_41(\uart_0|the_processor_uart_0_regs|readdata[4]~q ),
	.readdata_42(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[4]~q ),
	.av_readdata_4(\jtag_uart_0|av_readdata[4]~3_combout ),
	.av_readdata_3(\jtag_uart_0|av_readdata[3]~4_combout ),
	.src_payload24(\mm_interconnect_0|cmd_mux_002|src_payload~8_combout ),
	.readdata_31(\uart_0|the_processor_uart_0_regs|readdata[3]~q ),
	.readdata_32(\seg|readdata[3]~combout ),
	.av_readdata_2(\jtag_uart_0|av_readdata[2]~5_combout ),
	.readdata_21(\seg|readdata[2]~combout ),
	.src_payload25(\mm_interconnect_0|cmd_mux_002|src_payload~9_combout ),
	.readdata_27(\seg_en|readdata[2]~combout ),
	.readdata_28(\uart_0|the_processor_uart_0_regs|readdata[2]~q ),
	.src_payload26(\mm_interconnect_0|cmd_mux_002|src_payload~10_combout ),
	.readdata_5(\seg|readdata[5]~combout ),
	.readdata_51(\uart_0|the_processor_uart_0_regs|readdata[5]~q ),
	.readdata_52(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[5]~q ),
	.av_readdata_5(\jtag_uart_0|av_readdata[5]~6_combout ),
	.d_writedata_14(\nios2_gen2_0|cpu|d_writedata[14]~q ),
	.src_payload27(\mm_interconnect_0|cmd_mux_002|src_payload~11_combout ),
	.d_byteenable_1(\nios2_gen2_0|cpu|d_byteenable[1]~q ),
	.src_data_33(\mm_interconnect_0|cmd_mux_002|src_data[33]~combout ),
	.readdata_141(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[14]~q ),
	.woverflow(\jtag_uart_0|woverflow~q ),
	.d_writedata_15(\nios2_gen2_0|cpu|d_writedata[15]~q ),
	.src_payload28(\mm_interconnect_0|cmd_mux_002|src_payload~12_combout ),
	.readdata_15(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[15]~q ),
	.rvalid(\jtag_uart_0|rvalid~q ),
	.d_writedata_11(\nios2_gen2_0|cpu|d_writedata[11]~q ),
	.src_payload29(\mm_interconnect_0|cmd_mux_002|src_payload~13_combout ),
	.readdata_111(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[11]~q ),
	.d_writedata_13(\nios2_gen2_0|cpu|d_writedata[13]~q ),
	.src_payload30(\mm_interconnect_0|cmd_mux_002|src_payload~14_combout ),
	.readdata_131(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[13]~q ),
	.d_writedata_16(\nios2_gen2_0|cpu|d_writedata[16]~q ),
	.src_payload31(\mm_interconnect_0|cmd_mux_002|src_payload~15_combout ),
	.readdata_16(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[16]~q ),
	.counter_reg_bit_01(\jtag_uart_0|the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.d_writedata_12(\nios2_gen2_0|cpu|d_writedata[12]~q ),
	.src_payload32(\mm_interconnect_0|cmd_mux_002|src_payload~16_combout ),
	.readdata_121(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[12]~q ),
	.b_non_empty(\jtag_uart_0|the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.av_readdata_pre_271(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[27]~q ),
	.av_readdata_pre_281(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[28]~q ),
	.av_readdata_pre_291(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[29]~q ),
	.av_readdata_pre_30(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[30]~q ),
	.av_readdata_pre_311(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[31]~q ),
	.d_writedata_10(\nios2_gen2_0|cpu|d_writedata[10]~q ),
	.src_payload33(\mm_interconnect_0|cmd_mux_002|src_payload~17_combout ),
	.readdata_10(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[10]~q ),
	.ac(\jtag_uart_0|ac~q ),
	.readdata_9(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[9]~q ),
	.readdata_91(\uart_0|the_processor_uart_0_regs|readdata[9]~q ),
	.src_payload34(\mm_interconnect_0|cmd_mux_002|src_payload~18_combout ),
	.readdata_8(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[8]~q ),
	.readdata_81(\uart_0|the_processor_uart_0_regs|readdata[8]~q ),
	.d_writedata_8(\nios2_gen2_0|cpu|d_writedata[8]~q ),
	.src_payload35(\mm_interconnect_0|cmd_mux_002|src_payload~19_combout ),
	.readdata_7(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[7]~q ),
	.av_readdata_7(\jtag_uart_0|av_readdata[7]~7_combout ),
	.src_payload36(\mm_interconnect_0|cmd_mux_002|src_payload~20_combout ),
	.readdata_71(\seg|readdata[7]~combout ),
	.readdata_72(\uart_0|the_processor_uart_0_regs|readdata[7]~q ),
	.readdata_6(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[6]~q ),
	.av_readdata_6(\jtag_uart_0|av_readdata[6]~8_combout ),
	.src_payload37(\mm_interconnect_0|cmd_mux_002|src_payload~21_combout ),
	.readdata_61(\seg|readdata[6]~combout ),
	.readdata_62(\uart_0|the_processor_uart_0_regs|readdata[6]~q ),
	.src_payload38(\mm_interconnect_0|rsp_mux|src_payload~2_combout ),
	.d_writedata_21(\nios2_gen2_0|cpu|d_writedata[21]~q ),
	.src_payload39(\mm_interconnect_0|cmd_mux_002|src_payload~22_combout ),
	.readdata_211(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[21]~q ),
	.counter_reg_bit_51(\jtag_uart_0|the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.d_writedata_20(\nios2_gen2_0|cpu|d_writedata[20]~q ),
	.src_payload40(\mm_interconnect_0|cmd_mux_002|src_payload~23_combout ),
	.readdata_20(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[20]~q ),
	.counter_reg_bit_41(\jtag_uart_0|the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.src_payload41(\mm_interconnect_0|rsp_mux|src_payload~4_combout ),
	.d_writedata_19(\nios2_gen2_0|cpu|d_writedata[19]~q ),
	.src_payload42(\mm_interconnect_0|cmd_mux_002|src_payload~24_combout ),
	.readdata_19(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[19]~q ),
	.counter_reg_bit_31(\jtag_uart_0|the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.src_payload43(\mm_interconnect_0|rsp_mux|src_payload~6_combout ),
	.d_writedata_18(\nios2_gen2_0|cpu|d_writedata[18]~q ),
	.src_payload44(\mm_interconnect_0|cmd_mux_002|src_payload~25_combout ),
	.counter_reg_bit_21(\jtag_uart_0|the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.readdata_18(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[18]~q ),
	.src_payload45(\mm_interconnect_0|rsp_mux|src_payload~8_combout ),
	.d_writedata_17(\nios2_gen2_0|cpu|d_writedata[17]~q ),
	.src_payload46(\mm_interconnect_0|cmd_mux_002|src_payload~26_combout ),
	.counter_reg_bit_11(\jtag_uart_0|the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.readdata_17(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[17]~q ),
	.src_payload47(\mm_interconnect_0|rsp_mux|src_payload~10_combout ),
	.src_payload48(\mm_interconnect_0|rsp_mux|src_payload~11_combout ),
	.src_payload49(\mm_interconnect_0|rsp_mux|src_payload~13_combout ),
	.src_data_9(\mm_interconnect_0|rsp_mux|src_data[9]~8_combout ),
	.end_begintransfer(\mm_interconnect_0|uart_0_s1_translator|end_begintransfer~q ),
	.src_data_382(\mm_interconnect_0|cmd_mux|src_data[38]~combout ),
	.src_payload50(\mm_interconnect_0|cmd_mux|src_payload~0_combout ),
	.src_payload51(\mm_interconnect_0|cmd_mux_001|src_payload~0_combout ),
	.src_payload52(\mm_interconnect_0|cmd_mux_001|src_payload~1_combout ),
	.src_data_383(\mm_interconnect_0|cmd_mux_001|src_data[38]~combout ),
	.src_data_392(\mm_interconnect_0|cmd_mux_001|src_data[39]~combout ),
	.src_data_402(\mm_interconnect_0|cmd_mux_001|src_data[40]~combout ),
	.src_data_411(\mm_interconnect_0|cmd_mux_001|src_data[41]~combout ),
	.src_data_421(\mm_interconnect_0|cmd_mux_001|src_data[42]~combout ),
	.src_data_431(\mm_interconnect_0|cmd_mux_001|src_data[43]~combout ),
	.src_data_441(\mm_interconnect_0|cmd_mux_001|src_data[44]~combout ),
	.src_data_451(\mm_interconnect_0|cmd_mux_001|src_data[45]~combout ),
	.src_data_321(\mm_interconnect_0|cmd_mux_001|src_data[32]~combout ),
	.src_payload53(\mm_interconnect_0|cmd_mux|src_payload~1_combout ),
	.src_payload54(\mm_interconnect_0|cmd_mux|src_payload~2_combout ),
	.readdata_271(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[27]~q ),
	.src_payload55(\mm_interconnect_0|cmd_mux_002|src_payload~27_combout ),
	.readdata_281(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[28]~q ),
	.src_payload56(\mm_interconnect_0|cmd_mux_002|src_payload~28_combout ),
	.readdata_29(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[29]~q ),
	.src_payload57(\mm_interconnect_0|cmd_mux_002|src_payload~29_combout ),
	.readdata_30(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[30]~q ),
	.src_payload58(\mm_interconnect_0|cmd_mux_002|src_payload~30_combout ),
	.readdata_311(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|readdata[31]~q ),
	.src_payload59(\mm_interconnect_0|cmd_mux_002|src_payload~31_combout ),
	.src_payload60(\mm_interconnect_0|rsp_mux|src_payload~14_combout ),
	.src_payload61(\mm_interconnect_0|rsp_mux|src_payload~16_combout ),
	.src_payload62(\mm_interconnect_0|rsp_mux|src_payload~18_combout ),
	.src_payload63(\mm_interconnect_0|rsp_mux|src_payload~20_combout ),
	.src_payload64(\mm_interconnect_0|rsp_mux|src_payload~22_combout ),
	.src_payload65(\mm_interconnect_0|rsp_mux|src_payload~24_combout ),
	.src_payload66(\mm_interconnect_0|rsp_mux|src_payload~26_combout ),
	.src_payload67(\mm_interconnect_0|cmd_mux_001|src_payload~2_combout ),
	.src_payload68(\mm_interconnect_0|cmd_mux_007|src_payload~9_combout ),
	.src_payload69(\mm_interconnect_0|cmd_mux_001|src_payload~3_combout ),
	.src_payload70(\mm_interconnect_0|cmd_mux_001|src_payload~4_combout ),
	.src_payload71(\mm_interconnect_0|cmd_mux_001|src_payload~5_combout ),
	.src_data_341(\mm_interconnect_0|cmd_mux_001|src_data[34]~combout ),
	.src_payload72(\mm_interconnect_0|cmd_mux_001|src_payload~6_combout ),
	.src_payload73(\mm_interconnect_0|cmd_mux_001|src_payload~7_combout ),
	.src_data_351(\mm_interconnect_0|cmd_mux_001|src_data[35]~combout ),
	.src_payload74(\mm_interconnect_0|cmd_mux_001|src_payload~8_combout ),
	.src_payload75(\mm_interconnect_0|cmd_mux_001|src_payload~9_combout ),
	.src_payload76(\mm_interconnect_0|cmd_mux_001|src_payload~10_combout ),
	.src_payload77(\mm_interconnect_0|cmd_mux_001|src_payload~11_combout ),
	.src_payload78(\mm_interconnect_0|cmd_mux_001|src_payload~12_combout ),
	.src_data_331(\mm_interconnect_0|cmd_mux_001|src_data[33]~combout ),
	.src_payload79(\mm_interconnect_0|cmd_mux_001|src_payload~13_combout ),
	.src_payload80(\mm_interconnect_0|cmd_mux_001|src_payload~14_combout ),
	.src_payload81(\mm_interconnect_0|cmd_mux_001|src_payload~15_combout ),
	.src_payload82(\mm_interconnect_0|cmd_mux_001|src_payload~16_combout ),
	.src_payload83(\mm_interconnect_0|cmd_mux_001|src_payload~17_combout ),
	.src_payload84(\mm_interconnect_0|cmd_mux_001|src_payload~18_combout ),
	.src_payload85(\mm_interconnect_0|cmd_mux_001|src_payload~19_combout ),
	.src_payload86(\mm_interconnect_0|cmd_mux_001|src_payload~20_combout ),
	.src_payload87(\mm_interconnect_0|cmd_mux_001|src_payload~21_combout ),
	.src_payload88(\mm_interconnect_0|cmd_mux_001|src_payload~22_combout ),
	.src_payload89(\mm_interconnect_0|cmd_mux_001|src_payload~23_combout ),
	.src_payload90(\mm_interconnect_0|cmd_mux_001|src_payload~24_combout ),
	.src_payload91(\mm_interconnect_0|cmd_mux_001|src_payload~25_combout ),
	.src_payload92(\mm_interconnect_0|cmd_mux_001|src_payload~26_combout ),
	.src_payload93(\mm_interconnect_0|cmd_mux_001|src_payload~27_combout ),
	.src_payload94(\mm_interconnect_0|cmd_mux|src_payload~3_combout ),
	.src_payload95(\mm_interconnect_0|cmd_mux_001|src_payload~28_combout ),
	.src_payload96(\mm_interconnect_0|cmd_mux_001|src_payload~29_combout ),
	.src_payload97(\mm_interconnect_0|cmd_mux_001|src_payload~30_combout ),
	.src_payload98(\mm_interconnect_0|cmd_mux_001|src_payload~31_combout ),
	.src_payload99(\mm_interconnect_0|cmd_mux_001|src_payload~32_combout ),
	.src_payload100(\mm_interconnect_0|cmd_mux|src_payload~4_combout ),
	.src_payload101(\mm_interconnect_0|cmd_mux|src_payload~5_combout ),
	.src_payload102(\mm_interconnect_0|cmd_mux|src_payload~6_combout ),
	.src_payload103(\mm_interconnect_0|cmd_mux|src_payload~7_combout ),
	.clk_clk(\clk_clk~input_o ));

processor_processor_uart_0 uart_0(
	.txd(\uart_0|the_processor_uart_0_tx|txd~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.mem_used_1(\mm_interconnect_0|uart_0_s1_agent_rsp_fifo|mem_used[1]~q ),
	.wait_latency_counter_1(\mm_interconnect_0|uart_0_s1_translator|wait_latency_counter[1]~q ),
	.src_payload(\mm_interconnect_0|cmd_mux_007|src_payload~0_combout ),
	.src_data_38(\mm_interconnect_0|cmd_mux_007|src_data[38]~combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux_007|src_data[39]~combout ),
	.src_data_40(\mm_interconnect_0|cmd_mux_007|src_data[40]~combout ),
	.WideOr1(\mm_interconnect_0|cmd_mux_007|WideOr1~combout ),
	.av_begintransfer(\mm_interconnect_0|uart_0_s1_translator|av_begintransfer~0_combout ),
	.src_data_56(\mm_interconnect_0|cmd_mux_007|src_data[56]~combout ),
	.rx_rd_strobe_onset(\uart_0|the_processor_uart_0_rx|rx_rd_strobe_onset~0_combout ),
	.src_payload1(\mm_interconnect_0|cmd_mux_007|src_payload~1_combout ),
	.src_payload2(\mm_interconnect_0|cmd_mux_007|src_payload~2_combout ),
	.src_payload3(\mm_interconnect_0|cmd_mux_007|src_payload~3_combout ),
	.src_payload4(\mm_interconnect_0|cmd_mux_007|src_payload~4_combout ),
	.src_payload5(\mm_interconnect_0|cmd_mux_007|src_payload~5_combout ),
	.src_payload6(\mm_interconnect_0|cmd_mux_007|src_payload~6_combout ),
	.src_payload7(\mm_interconnect_0|cmd_mux_007|src_payload~7_combout ),
	.src_payload8(\mm_interconnect_0|cmd_mux_007|src_payload~8_combout ),
	.readdata_0(\uart_0|the_processor_uart_0_regs|readdata[0]~q ),
	.irq(\uart_0|the_processor_uart_0_regs|irq~q ),
	.readdata_1(\uart_0|the_processor_uart_0_regs|readdata[1]~q ),
	.readdata_4(\uart_0|the_processor_uart_0_regs|readdata[4]~q ),
	.readdata_3(\uart_0|the_processor_uart_0_regs|readdata[3]~q ),
	.readdata_2(\uart_0|the_processor_uart_0_regs|readdata[2]~q ),
	.readdata_5(\uart_0|the_processor_uart_0_regs|readdata[5]~q ),
	.readdata_9(\uart_0|the_processor_uart_0_regs|readdata[9]~q ),
	.readdata_8(\uart_0|the_processor_uart_0_regs|readdata[8]~q ),
	.readdata_7(\uart_0|the_processor_uart_0_regs|readdata[7]~q ),
	.readdata_6(\uart_0|the_processor_uart_0_regs|readdata[6]~q ),
	.end_begintransfer(\mm_interconnect_0|uart_0_s1_translator|end_begintransfer~q ),
	.src_payload9(\mm_interconnect_0|cmd_mux_007|src_payload~9_combout ),
	.GND_port(\~GND~combout ),
	.clk_clk(\clk_clk~input_o ),
	.uart_0_rxd(\uart_0_rxd~input_o ));

processor_processor_onchip_memory2_0 onchip_memory2_0(
	.q_a_0(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[0] ),
	.q_a_22(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_23(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_24(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[24] ),
	.q_a_25(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[25] ),
	.q_a_26(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[26] ),
	.q_a_1(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[1] ),
	.q_a_4(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[4] ),
	.q_a_3(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[3] ),
	.q_a_2(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[2] ),
	.q_a_5(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_14(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_15(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_11(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_13(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_16(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[16] ),
	.q_a_12(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_10(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_9(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_8(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_7(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[7] ),
	.q_a_6(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[6] ),
	.q_a_21(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[21] ),
	.q_a_20(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[20] ),
	.q_a_19(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[19] ),
	.q_a_18(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[18] ),
	.q_a_17(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[17] ),
	.q_a_27(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[27] ),
	.q_a_28(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[28] ),
	.q_a_29(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[29] ),
	.q_a_30(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[30] ),
	.q_a_31(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[31] ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_002|saved_grant[0]~q ),
	.mem_used_1(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem_used[1]~q ),
	.uav_write(\mm_interconnect_0|nios2_gen2_0_data_master_translator|uav_write~0_combout ),
	.WideOr1(\mm_interconnect_0|cmd_mux_002|WideOr1~combout ),
	.r_early_rst(\rst_controller|r_early_rst~q ),
	.src_payload(\mm_interconnect_0|cmd_mux_002|src_payload~0_combout ),
	.src_data_38(\mm_interconnect_0|cmd_mux_002|src_data[38]~combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux_002|src_data[39]~combout ),
	.src_data_40(\mm_interconnect_0|cmd_mux_002|src_data[40]~combout ),
	.src_data_41(\mm_interconnect_0|cmd_mux_002|src_data[41]~combout ),
	.src_data_42(\mm_interconnect_0|cmd_mux_002|src_data[42]~combout ),
	.src_data_43(\mm_interconnect_0|cmd_mux_002|src_data[43]~combout ),
	.src_data_44(\mm_interconnect_0|cmd_mux_002|src_data[44]~combout ),
	.src_data_45(\mm_interconnect_0|cmd_mux_002|src_data[45]~combout ),
	.src_data_46(\mm_interconnect_0|cmd_mux_002|src_data[46]~combout ),
	.src_data_47(\mm_interconnect_0|cmd_mux_002|src_data[47]~combout ),
	.src_data_48(\mm_interconnect_0|cmd_mux_002|src_data[48]~combout ),
	.src_data_49(\mm_interconnect_0|cmd_mux_002|src_data[49]~combout ),
	.src_data_50(\mm_interconnect_0|cmd_mux_002|src_data[50]~combout ),
	.src_data_32(\mm_interconnect_0|cmd_mux_002|src_data[32]~combout ),
	.src_payload1(\mm_interconnect_0|cmd_mux_002|src_payload~1_combout ),
	.src_data_34(\mm_interconnect_0|cmd_mux_002|src_data[34]~combout ),
	.src_payload2(\mm_interconnect_0|cmd_mux_002|src_payload~2_combout ),
	.src_payload3(\mm_interconnect_0|cmd_mux_002|src_payload~3_combout ),
	.src_data_35(\mm_interconnect_0|cmd_mux_002|src_data[35]~combout ),
	.src_payload4(\mm_interconnect_0|cmd_mux_002|src_payload~4_combout ),
	.src_payload5(\mm_interconnect_0|cmd_mux_002|src_payload~5_combout ),
	.src_payload6(\mm_interconnect_0|cmd_mux_002|src_payload~6_combout ),
	.src_payload7(\mm_interconnect_0|cmd_mux_002|src_payload~7_combout ),
	.src_payload8(\mm_interconnect_0|cmd_mux_002|src_payload~8_combout ),
	.src_payload9(\mm_interconnect_0|cmd_mux_002|src_payload~9_combout ),
	.src_payload10(\mm_interconnect_0|cmd_mux_002|src_payload~10_combout ),
	.src_payload11(\mm_interconnect_0|cmd_mux_002|src_payload~11_combout ),
	.src_data_33(\mm_interconnect_0|cmd_mux_002|src_data[33]~combout ),
	.src_payload12(\mm_interconnect_0|cmd_mux_002|src_payload~12_combout ),
	.src_payload13(\mm_interconnect_0|cmd_mux_002|src_payload~13_combout ),
	.src_payload14(\mm_interconnect_0|cmd_mux_002|src_payload~14_combout ),
	.src_payload15(\mm_interconnect_0|cmd_mux_002|src_payload~15_combout ),
	.src_payload16(\mm_interconnect_0|cmd_mux_002|src_payload~16_combout ),
	.src_payload17(\mm_interconnect_0|cmd_mux_002|src_payload~17_combout ),
	.src_payload18(\mm_interconnect_0|cmd_mux_002|src_payload~18_combout ),
	.src_payload19(\mm_interconnect_0|cmd_mux_002|src_payload~19_combout ),
	.src_payload20(\mm_interconnect_0|cmd_mux_002|src_payload~20_combout ),
	.src_payload21(\mm_interconnect_0|cmd_mux_002|src_payload~21_combout ),
	.src_payload22(\mm_interconnect_0|cmd_mux_002|src_payload~22_combout ),
	.src_payload23(\mm_interconnect_0|cmd_mux_002|src_payload~23_combout ),
	.src_payload24(\mm_interconnect_0|cmd_mux_002|src_payload~24_combout ),
	.src_payload25(\mm_interconnect_0|cmd_mux_002|src_payload~25_combout ),
	.src_payload26(\mm_interconnect_0|cmd_mux_002|src_payload~26_combout ),
	.src_payload27(\mm_interconnect_0|cmd_mux_002|src_payload~27_combout ),
	.src_payload28(\mm_interconnect_0|cmd_mux_002|src_payload~28_combout ),
	.src_payload29(\mm_interconnect_0|cmd_mux_002|src_payload~29_combout ),
	.src_payload30(\mm_interconnect_0|cmd_mux_002|src_payload~30_combout ),
	.src_payload31(\mm_interconnect_0|cmd_mux_002|src_payload~31_combout ),
	.clk_clk(\clk_clk~input_o ));

processor_altera_reset_controller rst_controller(
	.r_sync_rst1(\rst_controller|r_sync_rst~q ),
	.r_early_rst1(\rst_controller|r_early_rst~q ),
	.altera_reset_synchronizer_int_chain_1(\rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ),
	.clk_clk(\clk_clk~input_o ),
	.reset_reset_n(\reset_reset_n~input_o ));

processor_processor_jtag_uart_0 jtag_uart_0(
	.adapted_tdo(\jtag_uart_0|processor_jtag_uart_0_alt_jtag_atlantic|adapted_tdo~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.rst1(\jtag_uart_0|processor_jtag_uart_0_alt_jtag_atlantic|rst1~q ),
	.av_waitrequest1(\jtag_uart_0|av_waitrequest~q ),
	.mem_used_1(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo|mem_used[1]~q ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux|saved_grant[0]~q ),
	.uav_write(\mm_interconnect_0|nios2_gen2_0_data_master_translator|uav_write~0_combout ),
	.src_data_56(\mm_interconnect_0|cmd_mux|src_data[56]~combout ),
	.WideOr1(\mm_interconnect_0|cmd_mux|WideOr1~combout ),
	.b_full(\jtag_uart_0|the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.read_01(\jtag_uart_0|read_0~q ),
	.av_readdata_0(\jtag_uart_0|av_readdata[0]~0_combout ),
	.av_readdata_9(\jtag_uart_0|av_readdata[9]~combout ),
	.av_readdata_8(\jtag_uart_0|av_readdata[8]~1_combout ),
	.b_full1(\jtag_uart_0|the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.counter_reg_bit_5(\jtag_uart_0|the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.counter_reg_bit_4(\jtag_uart_0|the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\jtag_uart_0|the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\jtag_uart_0|the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\jtag_uart_0|the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\jtag_uart_0|the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.av_readdata_1(\jtag_uart_0|av_readdata[1]~2_combout ),
	.av_readdata_4(\jtag_uart_0|av_readdata[4]~3_combout ),
	.av_readdata_3(\jtag_uart_0|av_readdata[3]~4_combout ),
	.av_readdata_2(\jtag_uart_0|av_readdata[2]~5_combout ),
	.av_readdata_5(\jtag_uart_0|av_readdata[5]~6_combout ),
	.woverflow1(\jtag_uart_0|woverflow~q ),
	.rvalid1(\jtag_uart_0|rvalid~q ),
	.counter_reg_bit_01(\jtag_uart_0|the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.b_non_empty(\jtag_uart_0|the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.d_writedata_10(\nios2_gen2_0|cpu|d_writedata[10]~q ),
	.ac1(\jtag_uart_0|ac~q ),
	.av_readdata_7(\jtag_uart_0|av_readdata[7]~7_combout ),
	.av_readdata_6(\jtag_uart_0|av_readdata[6]~8_combout ),
	.counter_reg_bit_51(\jtag_uart_0|the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.counter_reg_bit_41(\jtag_uart_0|the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.counter_reg_bit_31(\jtag_uart_0|the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_21(\jtag_uart_0|the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.counter_reg_bit_11(\jtag_uart_0|the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.src_data_38(\mm_interconnect_0|cmd_mux|src_data[38]~combout ),
	.src_payload(\mm_interconnect_0|cmd_mux|src_payload~0_combout ),
	.src_payload1(\mm_interconnect_0|cmd_mux|src_payload~1_combout ),
	.src_payload2(\mm_interconnect_0|cmd_mux|src_payload~2_combout ),
	.src_payload3(\mm_interconnect_0|cmd_mux|src_payload~3_combout ),
	.src_payload4(\mm_interconnect_0|cmd_mux|src_payload~4_combout ),
	.src_payload5(\mm_interconnect_0|cmd_mux|src_payload~5_combout ),
	.src_payload6(\mm_interconnect_0|cmd_mux|src_payload~6_combout ),
	.src_payload7(\mm_interconnect_0|cmd_mux|src_payload~7_combout ),
	.altera_internal_jtag(\altera_internal_jtag~TCKUTAP ),
	.altera_internal_jtag1(\altera_internal_jtag~TDIUTAP ),
	.state_4(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.splitter_nodes_receive_0_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.virtual_ir_scan_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.clr_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.state_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.state_8(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.irf_reg_0_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.clk_clk(\clk_clk~input_o ));

processor_processor_SW sw(
	.W_alu_result_2(\nios2_gen2_0|cpu|W_alu_result[2]~q ),
	.W_alu_result_3(\nios2_gen2_0|cpu|W_alu_result[3]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.F_pc_1(\nios2_gen2_0|cpu|F_pc[1]~q ),
	.F_pc_0(\nios2_gen2_0|cpu|F_pc[0]~q ),
	.read_mux_out(\sw|read_mux_out~0_combout ),
	.read_mux_out1(\sw|read_mux_out~1_combout ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_006|saved_grant[0]~q ),
	.saved_grant_1(\mm_interconnect_0|cmd_mux_006|saved_grant[1]~q ),
	.readdata_0(\sw|readdata[0]~q ),
	.clk_clk(\clk_clk~input_o ),
	.sw_export(\sw_export~input_o ));

processor_processor_SEG_EN seg_en(
	.data_out_0(\seg_en|data_out[0]~q ),
	.data_out_1(\seg_en|data_out[1]~q ),
	.data_out_2(\seg_en|data_out[2]~q ),
	.writedata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\nios2_gen2_0|cpu|d_writedata[2]~q ,\nios2_gen2_0|cpu|d_writedata[1]~q ,\nios2_gen2_0|cpu|d_writedata[0]~q }),
	.reset_n(\rst_controller|r_sync_rst~q ),
	.read_mux_out(\sw|read_mux_out~0_combout ),
	.read_mux_out1(\sw|read_mux_out~1_combout ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_004|saved_grant[0]~q ),
	.src_payload(\mm_interconnect_0|cmd_mux_004|src_payload~0_combout ),
	.saved_grant_1(\mm_interconnect_0|cmd_mux_004|saved_grant[1]~q ),
	.src_valid(\mm_interconnect_0|cmd_mux_004|src_valid~3_combout ),
	.src_valid1(\mm_interconnect_0|cmd_mux_004|src_valid~5_combout ),
	.mem_used_1(\mm_interconnect_0|seg_en_s1_agent_rsp_fifo|mem_used[1]~q ),
	.always0(\seg_en|always0~0_combout ),
	.wait_latency_counter_1(\mm_interconnect_0|seg_en_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|seg_en_s1_translator|wait_latency_counter[0]~q ),
	.readdata_0(\seg_en|readdata[0]~combout ),
	.readdata_1(\seg_en|readdata[1]~combout ),
	.readdata_2(\seg_en|readdata[2]~combout ),
	.clk(\clk_clk~input_o ));

processor_processor_SEG seg(
	.data_out_0(\seg|data_out[0]~q ),
	.data_out_1(\seg|data_out[1]~q ),
	.data_out_2(\seg|data_out[2]~q ),
	.data_out_3(\seg|data_out[3]~q ),
	.data_out_4(\seg|data_out[4]~q ),
	.data_out_5(\seg|data_out[5]~q ),
	.data_out_6(\seg|data_out[6]~q ),
	.data_out_7(\seg|data_out[7]~q ),
	.writedata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\nios2_gen2_0|cpu|d_writedata[7]~q ,\nios2_gen2_0|cpu|d_writedata[6]~q ,\nios2_gen2_0|cpu|d_writedata[5]~q ,\nios2_gen2_0|cpu|d_writedata[4]~q ,\nios2_gen2_0|cpu|d_writedata[3]~q ,
\nios2_gen2_0|cpu|d_writedata[2]~q ,\nios2_gen2_0|cpu|d_writedata[1]~q ,\nios2_gen2_0|cpu|d_writedata[0]~q }),
	.reset_n(\rst_controller|r_sync_rst~q ),
	.read_mux_out(\sw|read_mux_out~0_combout ),
	.read_mux_out1(\sw|read_mux_out~1_combout ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_005|saved_grant[0]~q ),
	.src_payload(\mm_interconnect_0|cmd_mux_005|src_payload~0_combout ),
	.saved_grant_1(\mm_interconnect_0|cmd_mux_005|saved_grant[1]~q ),
	.src_valid(\mm_interconnect_0|cmd_mux_005|src_valid~2_combout ),
	.src_valid1(\mm_interconnect_0|cmd_mux_005|src_valid~4_combout ),
	.mem_used_1(\mm_interconnect_0|seg_s1_agent_rsp_fifo|mem_used[1]~q ),
	.always0(\seg|always0~0_combout ),
	.wait_latency_counter_1(\mm_interconnect_0|seg_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|seg_s1_translator|wait_latency_counter[0]~q ),
	.readdata_0(\seg|readdata[0]~combout ),
	.readdata_1(\seg|readdata[1]~combout ),
	.readdata_4(\seg|readdata[4]~combout ),
	.readdata_3(\seg|readdata[3]~combout ),
	.readdata_2(\seg|readdata[2]~combout ),
	.readdata_5(\seg|readdata[5]~combout ),
	.readdata_7(\seg|readdata[7]~combout ),
	.readdata_6(\seg|readdata[6]~combout ),
	.clk(\clk_clk~input_o ));

processor_processor_LED led(
	.data_out_0(\led|data_out[0]~q ),
	.data_out_1(\led|data_out[1]~q ),
	.d_writedata_0(\nios2_gen2_0|cpu|d_writedata[0]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_003|saved_grant[0]~q ),
	.src_payload(\mm_interconnect_0|cmd_mux_003|src_payload~0_combout ),
	.saved_grant_1(\mm_interconnect_0|cmd_mux_003|saved_grant[1]~q ),
	.src_valid(\mm_interconnect_0|cmd_mux_003|src_valid~3_combout ),
	.src_valid1(\mm_interconnect_0|cmd_mux_003|src_valid~5_combout ),
	.mem_used_1(\mm_interconnect_0|led_s1_agent_rsp_fifo|mem_used[1]~q ),
	.always0(\led|always0~0_combout ),
	.read_mux_out(\sw|read_mux_out~0_combout ),
	.read_mux_out1(\sw|read_mux_out~1_combout ),
	.wait_latency_counter_1(\mm_interconnect_0|led_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|led_s1_translator|wait_latency_counter[0]~q ),
	.d_writedata_1(\nios2_gen2_0|cpu|d_writedata[1]~q ),
	.readdata_0(\led|readdata[0]~combout ),
	.readdata_1(\led|readdata[1]~combout ),
	.clk(\clk_clk~input_o ));

cyclone10lp_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\~GND~combout ),
	.cout());
defparam \~GND .lut_mask = 16'h0000;
defparam \~GND .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~7_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~9_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~10_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~9_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 (
	.dataa(gnd),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .lut_mask = 16'h3FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.datab(\altera_internal_jtag~TDIUTAP ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .lut_mask = 16'hFFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(\altera_internal_jtag~TDIUTAP ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~5 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~5_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~6 .lut_mask = 16'hFFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~6 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~7_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~7 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0 .lut_mask = 16'hEEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~8 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~8_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~1_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~9 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~9 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~8_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~7_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~10 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~1 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~1_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~7 .lut_mask = 16'hFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~8 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~8 .sum_lutc_input = "datac";

assign \clk_clk~input_o  = clk_clk;

assign \sw_export~input_o  = sw_export;

assign \reset_reset_n~input_o  = reset_reset_n;

assign \uart_0_rxd~input_o  = uart_0_rxd;

assign led_export[0] = ~ \led|data_out[0]~q ;

assign led_export[1] = ~ \led|data_out[1]~q ;

assign seg_export[0] = \seg|data_out[0]~q ;

assign seg_export[1] = \seg|data_out[1]~q ;

assign seg_export[2] = \seg|data_out[2]~q ;

assign seg_export[3] = \seg|data_out[3]~q ;

assign seg_export[4] = \seg|data_out[4]~q ;

assign seg_export[5] = \seg|data_out[5]~q ;

assign seg_export[6] = \seg|data_out[6]~q ;

assign seg_export[7] = \seg|data_out[7]~q ;

assign seg_en_export[0] = \seg_en|data_out[0]~q ;

assign seg_en_export[1] = \seg_en|data_out[1]~q ;

assign seg_en_export[2] = \seg_en|data_out[2]~q ;

assign uart_0_txd = ~ \uart_0|the_processor_uart_0_tx|txd~q ;

assign altera_reserved_tdo = \altera_internal_jtag~TDO ;

assign \altera_reserved_tms~input_o  = altera_reserved_tms;

assign \altera_reserved_tck~input_o  = altera_reserved_tck;

assign \altera_reserved_tdi~input_o  = altera_reserved_tdi;

cyclone10lp_jtag altera_internal_jtag(
	.tms(\altera_reserved_tms~input_o ),
	.tck(\altera_reserved_tck~input_o ),
	.tdi(\altera_reserved_tdi~input_o ),
	.tdoutap(gnd),
	.tdouser(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.tdo(\altera_internal_jtag~TDO ),
	.tmsutap(\altera_internal_jtag~TMSUTAP ),
	.tckutap(\altera_internal_jtag~TCKUTAP ),
	.tdiutap(\altera_internal_jtag~TDIUTAP ),
	.shiftuser(),
	.clkdruser(),
	.updateuser(),
	.runidleuser(),
	.usr1user());

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TMSUTAP ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .lut_mask = 16'h0FF0;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .lut_mask = 16'hC33C;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .lut_mask = 16'hFF7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TMSUTAP ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .lut_mask = 16'h7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .lut_mask = 16'hEEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(\rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ),
	.datad(\rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~6 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~7 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~4 .lut_mask = 16'hEEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~6_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~7_combout ),
	.datac(\altera_internal_jtag~TDIUTAP ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~4_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~14 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~14_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~14 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9 (
	.dataa(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_tck|ir_out[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9 .lut_mask = 16'hFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~16_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~7 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~7 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~7_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~10 .lut_mask = 16'hFFB8;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~16 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~10_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~16_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~16 .lut_mask = 16'hFFAC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~16 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~14_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~16_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~15 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~15_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~15 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~15 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~15_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~16_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~13 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~13 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~13_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~16_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 .lut_mask = 16'h3FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~8 .lut_mask = 16'hF7FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3 .lut_mask = 16'h8B8B;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~8_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~4 .lut_mask = 16'hB8FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~4 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~4_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~14_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~5 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~5 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~1 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~1_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 .lut_mask = 16'hFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~4 .lut_mask = 16'hFFAC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~5 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~4_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~5_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~6 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~6 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~11 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12 (
	.dataa(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_tck|ir_out[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~11_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~16_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~6 .lut_mask = 16'hFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~6 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~6_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~4_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 (
	.dataa(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(\jtag_uart_0|processor_jtag_uart_0_alt_jtag_atlantic|adapted_tdo~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .lut_mask = 16'hFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~6 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5 .lut_mask = 16'h55AA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .lut_mask = 16'h3FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~15 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~15_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~15 .lut_mask = 16'hFFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~16 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~16_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~16 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~16 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~15_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~16_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~6 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~7_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~8 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~7 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~7 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~15_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~16_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~8 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~9_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~10 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~9 .lut_mask = 16'h5AAF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~9 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~15_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~16_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~10 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~11_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~12 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~11 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~11 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~15_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~16_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~12 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~13 .lut_mask = 16'h5A5A;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~13 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~15_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~16_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .lut_mask = 16'hFF96;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .lut_mask = 16'hD8D8;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~7 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~7_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~8 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~8_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .lut_mask = 16'h6FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~7_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~8_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13 .lut_mask = 16'hD77D;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14 .lut_mask = 16'hDEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~8_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11 .lut_mask = 16'h8BFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~8_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .lut_mask = 16'h0FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena .lut_mask = 16'hFFFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3_combout ),
	.asdata(\altera_internal_jtag~TDIUTAP ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~12 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11 .lut_mask = 16'h55AA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~12 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~23 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~23_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~23 .lut_mask = 16'hFFFB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~23 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~17 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16 .lut_mask = 16'h5AAF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~17 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~19 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~19 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20 .lut_mask = 16'h5A5A;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~15 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~15_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~15 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~22 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~15_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~22_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~22 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~22 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .lut_mask = 16'h7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~19 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~19_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~19 .lut_mask = 16'hFF6F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10 .lut_mask = 16'hAFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12 (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12 .lut_mask = 16'h3FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .lut_mask = 16'h3FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~14 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~14_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~14 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~15 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~15_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~15 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~17 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~17_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~17 .lut_mask = 16'hFFBF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~18 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~17_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~18_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~18 .lut_mask = 16'hBF8F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~16 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~14_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~15_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~16_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~16 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~16 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~19_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .lut_mask = 16'hFFBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .lut_mask = 16'hFFDF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1] .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 (
	.dataa(\jtag_uart_0|processor_jtag_uart_0_alt_jtag_atlantic|adapted_tdo~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .lut_mask = 16'hACFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ),
	.datab(\nios2_gen2_0|cpu|the_processor_nios2_gen2_0_cpu_nios2_oci|the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8 .lut_mask = 16'hAFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo (
	.clk(!\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .power_up = "low";

cyclone10lp_lcell_comb \auto_hub|~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|~GND~combout ),
	.cout());
defparam \auto_hub|~GND .lut_mask = 16'h0000;
defparam \auto_hub|~GND .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .sum_lutc_input = "datac";

endmodule

module processor_altera_reset_controller (
	r_sync_rst1,
	r_early_rst1,
	altera_reset_synchronizer_int_chain_1,
	clk_clk,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
output 	r_sync_rst1;
output 	r_early_rst1;
output 	altera_reset_synchronizer_int_chain_1;
input 	clk_clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;
wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[2]~q ;
wire \altera_reset_synchronizer_int_chain[3]~q ;
wire \altera_reset_synchronizer_int_chain[4]~0_combout ;
wire \altera_reset_synchronizer_int_chain[4]~q ;
wire \r_sync_rst_chain[3]~q ;
wire \r_sync_rst_chain~1_combout ;
wire \r_sync_rst_chain[2]~q ;
wire \r_sync_rst_chain~0_combout ;
wire \r_sync_rst_chain[1]~q ;
wire \WideOr0~0_combout ;
wire \always2~0_combout ;


processor_altera_reset_synchronizer alt_rst_req_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.altera_reset_synchronizer_int_chain_1(altera_reset_synchronizer_int_chain_1),
	.clk(clk_clk));

processor_altera_reset_synchronizer_1 alt_rst_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.clk(clk_clk),
	.reset_reset_n(reset_reset_n));

dffeas r_sync_rst(
	.clk(clk_clk),
	.d(\WideOr0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_sync_rst1),
	.prn(vcc));
defparam r_sync_rst.is_wysiwyg = "true";
defparam r_sync_rst.power_up = "low";

dffeas r_early_rst(
	.clk(clk_clk),
	.d(\always2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_early_rst1),
	.prn(vcc));
defparam r_early_rst.is_wysiwyg = "true";
defparam r_early_rst.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk_clk),
	.d(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[2] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[2]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[2] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[2] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[3] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[3]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[3] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[3] .power_up = "low";

cyclone10lp_lcell_comb \altera_reset_synchronizer_int_chain[4]~0 (
	.dataa(\altera_reset_synchronizer_int_chain[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.cout());
defparam \altera_reset_synchronizer_int_chain[4]~0 .lut_mask = 16'h5555;
defparam \altera_reset_synchronizer_int_chain[4]~0 .sum_lutc_input = "datac";

dffeas \altera_reset_synchronizer_int_chain[4] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[4]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[4] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[4] .power_up = "low";

dffeas \r_sync_rst_chain[3] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[3]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[3] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[3] .power_up = "low";

cyclone10lp_lcell_comb \r_sync_rst_chain~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_reset_synchronizer_int_chain[2]~q ),
	.datad(\r_sync_rst_chain[3]~q ),
	.cin(gnd),
	.combout(\r_sync_rst_chain~1_combout ),
	.cout());
defparam \r_sync_rst_chain~1 .lut_mask = 16'hFFF0;
defparam \r_sync_rst_chain~1 .sum_lutc_input = "datac";

dffeas \r_sync_rst_chain[2] (
	.clk(clk_clk),
	.d(\r_sync_rst_chain~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[2]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[2] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[2] .power_up = "low";

cyclone10lp_lcell_comb \r_sync_rst_chain~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_reset_synchronizer_int_chain[2]~q ),
	.datad(\r_sync_rst_chain[2]~q ),
	.cin(gnd),
	.combout(\r_sync_rst_chain~0_combout ),
	.cout());
defparam \r_sync_rst_chain~0 .lut_mask = 16'hFFF0;
defparam \r_sync_rst_chain~0 .sum_lutc_input = "datac";

dffeas \r_sync_rst_chain[1] (
	.clk(clk_clk),
	.d(\r_sync_rst_chain~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[1]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[1] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[1] .power_up = "low";

cyclone10lp_lcell_comb \WideOr0~0 (
	.dataa(\altera_reset_synchronizer_int_chain[4]~q ),
	.datab(r_sync_rst1),
	.datac(gnd),
	.datad(\r_sync_rst_chain[1]~q ),
	.cin(gnd),
	.combout(\WideOr0~0_combout ),
	.cout());
defparam \WideOr0~0 .lut_mask = 16'hEEFF;
defparam \WideOr0~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \always2~0 (
	.dataa(\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\r_sync_rst_chain[2]~q ),
	.cin(gnd),
	.combout(\always2~0_combout ),
	.cout());
defparam \always2~0 .lut_mask = 16'hAAFF;
defparam \always2~0 .sum_lutc_input = "datac";

endmodule

module processor_altera_reset_synchronizer (
	altera_reset_synchronizer_int_chain_out1,
	altera_reset_synchronizer_int_chain_1,
	clk)/* synthesis synthesis_greybox=1 */;
output 	altera_reset_synchronizer_int_chain_out1;
output 	altera_reset_synchronizer_int_chain_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

cyclone10lp_lcell_comb \altera_reset_synchronizer_int_chain[1]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(altera_reset_synchronizer_int_chain_1),
	.cout());
defparam \altera_reset_synchronizer_int_chain[1]~0 .lut_mask = 16'h0000;
defparam \altera_reset_synchronizer_int_chain[1]~0 .sum_lutc_input = "datac";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(altera_reset_synchronizer_int_chain_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module processor_altera_reset_synchronizer_1 (
	altera_reset_synchronizer_int_chain_out1,
	clk,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
output 	altera_reset_synchronizer_int_chain_out1;
input 	clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module processor_processor_jtag_uart_0 (
	adapted_tdo,
	r_sync_rst,
	rst1,
	av_waitrequest1,
	mem_used_1,
	saved_grant_0,
	uav_write,
	src_data_56,
	WideOr1,
	b_full,
	read_01,
	av_readdata_0,
	av_readdata_9,
	av_readdata_8,
	b_full1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	av_readdata_1,
	av_readdata_4,
	av_readdata_3,
	av_readdata_2,
	av_readdata_5,
	woverflow1,
	rvalid1,
	counter_reg_bit_01,
	b_non_empty,
	d_writedata_10,
	ac1,
	av_readdata_7,
	av_readdata_6,
	counter_reg_bit_51,
	counter_reg_bit_41,
	counter_reg_bit_31,
	counter_reg_bit_21,
	counter_reg_bit_11,
	src_data_38,
	src_payload,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	splitter_nodes_receive_0_3,
	virtual_ir_scan_reg,
	clr_reg,
	state_3,
	state_8,
	irf_reg_0_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	adapted_tdo;
input 	r_sync_rst;
output 	rst1;
output 	av_waitrequest1;
input 	mem_used_1;
input 	saved_grant_0;
input 	uav_write;
input 	src_data_56;
input 	WideOr1;
output 	b_full;
output 	read_01;
output 	av_readdata_0;
output 	av_readdata_9;
output 	av_readdata_8;
output 	b_full1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	av_readdata_1;
output 	av_readdata_4;
output 	av_readdata_3;
output 	av_readdata_2;
output 	av_readdata_5;
output 	woverflow1;
output 	rvalid1;
output 	counter_reg_bit_01;
output 	b_non_empty;
input 	d_writedata_10;
output 	ac1;
output 	av_readdata_7;
output 	av_readdata_6;
output 	counter_reg_bit_51;
output 	counter_reg_bit_41;
output 	counter_reg_bit_31;
output 	counter_reg_bit_21;
output 	counter_reg_bit_11;
input 	src_data_38;
input 	src_payload;
input 	src_payload1;
input 	src_payload2;
input 	src_payload3;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	splitter_nodes_receive_0_3;
input 	virtual_ir_scan_reg;
input 	clr_reg;
input 	state_3;
input 	state_8;
input 	irf_reg_0_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \t_dav~q ;
wire \processor_jtag_uart_0_alt_jtag_atlantic|rvalid0~q ;
wire \r_val~q ;
wire \processor_jtag_uart_0_alt_jtag_atlantic|r_ena1~q ;
wire \processor_jtag_uart_0_alt_jtag_atlantic|t_ena~reg0_q ;
wire \fifo_rd~1_combout ;
wire \the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ;
wire \r_val~0_combout ;
wire \fifo_wr~q ;
wire \wr_rfifo~combout ;
wire \processor_jtag_uart_0_alt_jtag_atlantic|wdata[0]~q ;
wire \processor_jtag_uart_0_alt_jtag_atlantic|t_pause~reg0_q ;
wire \processor_jtag_uart_0_alt_jtag_atlantic|wdata[1]~q ;
wire \processor_jtag_uart_0_alt_jtag_atlantic|wdata[4]~q ;
wire \processor_jtag_uart_0_alt_jtag_atlantic|wdata[3]~q ;
wire \processor_jtag_uart_0_alt_jtag_atlantic|wdata[2]~q ;
wire \processor_jtag_uart_0_alt_jtag_atlantic|wdata[5]~q ;
wire \processor_jtag_uart_0_alt_jtag_atlantic|wdata[7]~q ;
wire \processor_jtag_uart_0_alt_jtag_atlantic|wdata[6]~q ;
wire \fifo_wr~0_combout ;
wire \fifo_rd~0_combout ;
wire \av_waitrequest~0_combout ;
wire \fifo_rd~2_combout ;
wire \ien_AE~0_combout ;
wire \ien_AF~q ;
wire \LessThan0~0_combout ;
wire \LessThan0~1_combout ;
wire \fifo_AE~q ;
wire \ien_AE~q ;
wire \pause_irq~0_combout ;
wire \pause_irq~q ;
wire \Add0~1 ;
wire \Add0~3 ;
wire \Add0~4_combout ;
wire \Add0~0_combout ;
wire \Add0~2_combout ;
wire \LessThan1~0_combout ;
wire \Add0~5 ;
wire \Add0~6_combout ;
wire \Add0~7 ;
wire \Add0~8_combout ;
wire \LessThan1~1_combout ;
wire \Add0~9 ;
wire \Add0~10_combout ;
wire \Add0~11 ;
wire \Add0~12_combout ;
wire \LessThan1~2_combout ;
wire \fifo_AF~q ;
wire \woverflow~0_combout ;
wire \woverflow~1_combout ;
wire \rvalid~0_combout ;
wire \ac~0_combout ;
wire \ac~1_combout ;


processor_alt_jtag_atlantic processor_jtag_uart_0_alt_jtag_atlantic(
	.r_dat({\the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[7] ,\the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[6] ,\the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[5] ,
\the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[4] ,\the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[3] ,\the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[2] ,
\the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[1] ,\the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[0] }),
	.adapted_tdo1(adapted_tdo),
	.rst_n(r_sync_rst),
	.rst11(rst1),
	.t_dav(\t_dav~q ),
	.rvalid01(\processor_jtag_uart_0_alt_jtag_atlantic|rvalid0~q ),
	.r_val(\r_val~q ),
	.r_ena11(\processor_jtag_uart_0_alt_jtag_atlantic|r_ena1~q ),
	.t_ena(\processor_jtag_uart_0_alt_jtag_atlantic|t_ena~reg0_q ),
	.wdata_0(\processor_jtag_uart_0_alt_jtag_atlantic|wdata[0]~q ),
	.t_pause(\processor_jtag_uart_0_alt_jtag_atlantic|t_pause~reg0_q ),
	.wdata_1(\processor_jtag_uart_0_alt_jtag_atlantic|wdata[1]~q ),
	.wdata_4(\processor_jtag_uart_0_alt_jtag_atlantic|wdata[4]~q ),
	.wdata_3(\processor_jtag_uart_0_alt_jtag_atlantic|wdata[3]~q ),
	.wdata_2(\processor_jtag_uart_0_alt_jtag_atlantic|wdata[2]~q ),
	.wdata_5(\processor_jtag_uart_0_alt_jtag_atlantic|wdata[5]~q ),
	.wdata_7(\processor_jtag_uart_0_alt_jtag_atlantic|wdata[7]~q ),
	.wdata_6(\processor_jtag_uart_0_alt_jtag_atlantic|wdata[6]~q ),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.splitter_nodes_receive_0_3(splitter_nodes_receive_0_3),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.clr_reg(clr_reg),
	.state_3(state_3),
	.state_8(state_8),
	.irf_reg_0_1(irf_reg_0_1),
	.clk(clk_clk));

processor_processor_jtag_uart_0_scfifo_r the_processor_jtag_uart_0_scfifo_r(
	.q_b_0(\the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.q_b_1(\the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_4(\the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_3(\the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_2(\the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_5(\the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_7(\the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.q_b_6(\the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.r_sync_rst(r_sync_rst),
	.b_full(b_full),
	.counter_reg_bit_0(counter_reg_bit_01),
	.b_non_empty(b_non_empty),
	.counter_reg_bit_5(counter_reg_bit_51),
	.counter_reg_bit_4(counter_reg_bit_41),
	.counter_reg_bit_3(counter_reg_bit_31),
	.counter_reg_bit_2(counter_reg_bit_21),
	.counter_reg_bit_1(counter_reg_bit_11),
	.t_ena(\processor_jtag_uart_0_alt_jtag_atlantic|t_ena~reg0_q ),
	.fifo_rd(\fifo_rd~1_combout ),
	.wr_rfifo(\wr_rfifo~combout ),
	.wdata_0(\processor_jtag_uart_0_alt_jtag_atlantic|wdata[0]~q ),
	.fifo_rd1(\fifo_rd~2_combout ),
	.wdata_1(\processor_jtag_uart_0_alt_jtag_atlantic|wdata[1]~q ),
	.wdata_4(\processor_jtag_uart_0_alt_jtag_atlantic|wdata[4]~q ),
	.wdata_3(\processor_jtag_uart_0_alt_jtag_atlantic|wdata[3]~q ),
	.wdata_2(\processor_jtag_uart_0_alt_jtag_atlantic|wdata[2]~q ),
	.wdata_5(\processor_jtag_uart_0_alt_jtag_atlantic|wdata[5]~q ),
	.wdata_7(\processor_jtag_uart_0_alt_jtag_atlantic|wdata[7]~q ),
	.wdata_6(\processor_jtag_uart_0_alt_jtag_atlantic|wdata[6]~q ),
	.clk_clk(clk_clk));

processor_processor_jtag_uart_0_scfifo_w the_processor_jtag_uart_0_scfifo_w(
	.q_b_7(\the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.q_b_0(\the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.q_b_1(\the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_2(\the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_3(\the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_6(\the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.q_b_5(\the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_4(\the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.r_sync_rst(r_sync_rst),
	.b_full(b_full1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.b_non_empty(\the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.r_val(\r_val~0_combout ),
	.fifo_wr(\fifo_wr~q ),
	.src_payload(src_payload),
	.src_payload1(src_payload1),
	.src_payload2(src_payload2),
	.src_payload3(src_payload3),
	.src_payload4(src_payload4),
	.src_payload5(src_payload5),
	.src_payload6(src_payload6),
	.src_payload7(src_payload7),
	.clk_clk(clk_clk));

dffeas t_dav(
	.clk(clk_clk),
	.d(b_full),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\t_dav~q ),
	.prn(vcc));
defparam t_dav.is_wysiwyg = "true";
defparam t_dav.power_up = "low";

dffeas r_val(
	.clk(clk_clk),
	.d(\r_val~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_val~q ),
	.prn(vcc));
defparam r_val.is_wysiwyg = "true";
defparam r_val.power_up = "low";

cyclone10lp_lcell_comb \fifo_rd~1 (
	.dataa(src_data_56),
	.datab(\fifo_rd~0_combout ),
	.datac(b_non_empty),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\fifo_rd~1_combout ),
	.cout());
defparam \fifo_rd~1 .lut_mask = 16'hFEFF;
defparam \fifo_rd~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \r_val~0 (
	.dataa(\the_processor_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.datab(\r_val~q ),
	.datac(\processor_jtag_uart_0_alt_jtag_atlantic|r_ena1~q ),
	.datad(\processor_jtag_uart_0_alt_jtag_atlantic|rvalid0~q ),
	.cin(gnd),
	.combout(\r_val~0_combout ),
	.cout());
defparam \r_val~0 .lut_mask = 16'hBFFF;
defparam \r_val~0 .sum_lutc_input = "datac";

dffeas fifo_wr(
	.clk(clk_clk),
	.d(\fifo_wr~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_wr~q ),
	.prn(vcc));
defparam fifo_wr.is_wysiwyg = "true";
defparam fifo_wr.power_up = "low";

cyclone10lp_lcell_comb wr_rfifo(
	.dataa(\processor_jtag_uart_0_alt_jtag_atlantic|t_ena~reg0_q ),
	.datab(gnd),
	.datac(gnd),
	.datad(b_full),
	.cin(gnd),
	.combout(\wr_rfifo~combout ),
	.cout());
defparam wr_rfifo.lut_mask = 16'hAAFF;
defparam wr_rfifo.sum_lutc_input = "datac";

cyclone10lp_lcell_comb \fifo_wr~0 (
	.dataa(b_full1),
	.datab(gnd),
	.datac(gnd),
	.datad(\woverflow~0_combout ),
	.cin(gnd),
	.combout(\fifo_wr~0_combout ),
	.cout());
defparam \fifo_wr~0 .lut_mask = 16'hFF55;
defparam \fifo_wr~0 .sum_lutc_input = "datac";

dffeas av_waitrequest(
	.clk(clk_clk),
	.d(\av_waitrequest~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_waitrequest1),
	.prn(vcc));
defparam av_waitrequest.is_wysiwyg = "true";
defparam av_waitrequest.power_up = "low";

dffeas read_0(
	.clk(clk_clk),
	.d(\fifo_rd~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_01),
	.prn(vcc));
defparam read_0.is_wysiwyg = "true";
defparam read_0.power_up = "low";

cyclone10lp_lcell_comb \av_readdata[0]~0 (
	.dataa(\the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.datab(\ien_AF~q ),
	.datac(gnd),
	.datad(read_01),
	.cin(gnd),
	.combout(av_readdata_0),
	.cout());
defparam \av_readdata[0]~0 .lut_mask = 16'hAACC;
defparam \av_readdata[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_readdata[9] (
	.dataa(\fifo_AE~q ),
	.datab(\ien_AE~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_9),
	.cout());
defparam \av_readdata[9] .lut_mask = 16'hEEEE;
defparam \av_readdata[9] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_readdata[8]~1 (
	.dataa(\ien_AF~q ),
	.datab(\pause_irq~q ),
	.datac(\fifo_AF~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_8),
	.cout());
defparam \av_readdata[8]~1 .lut_mask = 16'hFEFE;
defparam \av_readdata[8]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_readdata[1]~2 (
	.dataa(\the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.datab(\ien_AE~q ),
	.datac(gnd),
	.datad(read_01),
	.cin(gnd),
	.combout(av_readdata_1),
	.cout());
defparam \av_readdata[1]~2 .lut_mask = 16'hAACC;
defparam \av_readdata[1]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_readdata[4]~3 (
	.dataa(read_01),
	.datab(\the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_4),
	.cout());
defparam \av_readdata[4]~3 .lut_mask = 16'hEEEE;
defparam \av_readdata[4]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_readdata[3]~4 (
	.dataa(read_01),
	.datab(\the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_3),
	.cout());
defparam \av_readdata[3]~4 .lut_mask = 16'hEEEE;
defparam \av_readdata[3]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_readdata[2]~5 (
	.dataa(read_01),
	.datab(\the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_2),
	.cout());
defparam \av_readdata[2]~5 .lut_mask = 16'hEEEE;
defparam \av_readdata[2]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_readdata[5]~6 (
	.dataa(read_01),
	.datab(\the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_5),
	.cout());
defparam \av_readdata[5]~6 .lut_mask = 16'hEEEE;
defparam \av_readdata[5]~6 .sum_lutc_input = "datac";

dffeas woverflow(
	.clk(clk_clk),
	.d(\woverflow~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(woverflow1),
	.prn(vcc));
defparam woverflow.is_wysiwyg = "true";
defparam woverflow.power_up = "low";

dffeas rvalid(
	.clk(clk_clk),
	.d(\rvalid~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rvalid1),
	.prn(vcc));
defparam rvalid.is_wysiwyg = "true";
defparam rvalid.power_up = "low";

dffeas ac(
	.clk(clk_clk),
	.d(\ac~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ac1),
	.prn(vcc));
defparam ac.is_wysiwyg = "true";
defparam ac.power_up = "low";

cyclone10lp_lcell_comb \av_readdata[7]~7 (
	.dataa(read_01),
	.datab(\the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_7),
	.cout());
defparam \av_readdata[7]~7 .lut_mask = 16'hEEEE;
defparam \av_readdata[7]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_readdata[6]~8 (
	.dataa(read_01),
	.datab(\the_processor_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_6),
	.cout());
defparam \av_readdata[6]~8 .lut_mask = 16'hEEEE;
defparam \av_readdata[6]~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \fifo_rd~0 (
	.dataa(WideOr1),
	.datab(gnd),
	.datac(av_waitrequest1),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\fifo_rd~0_combout ),
	.cout());
defparam \fifo_rd~0 .lut_mask = 16'hAFFF;
defparam \fifo_rd~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_waitrequest~0 (
	.dataa(\fifo_rd~0_combout ),
	.datab(src_data_56),
	.datac(uav_write),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(\av_waitrequest~0_combout ),
	.cout());
defparam \av_waitrequest~0 .lut_mask = 16'hFFFE;
defparam \av_waitrequest~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \fifo_rd~2 (
	.dataa(src_data_56),
	.datab(\fifo_rd~0_combout ),
	.datac(gnd),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\fifo_rd~2_combout ),
	.cout());
defparam \fifo_rd~2 .lut_mask = 16'hEEFF;
defparam \fifo_rd~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ien_AE~0 (
	.dataa(uav_write),
	.datab(saved_grant_0),
	.datac(\fifo_rd~0_combout ),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\ien_AE~0_combout ),
	.cout());
defparam \ien_AE~0 .lut_mask = 16'hFFFE;
defparam \ien_AE~0 .sum_lutc_input = "datac";

dffeas ien_AF(
	.clk(clk_clk),
	.d(src_payload1),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ien_AE~0_combout ),
	.q(\ien_AF~q ),
	.prn(vcc));
defparam ien_AF.is_wysiwyg = "true";
defparam ien_AF.power_up = "low";

cyclone10lp_lcell_comb \LessThan0~0 (
	.dataa(counter_reg_bit_3),
	.datab(counter_reg_bit_2),
	.datac(counter_reg_bit_1),
	.datad(counter_reg_bit_0),
	.cin(gnd),
	.combout(\LessThan0~0_combout ),
	.cout());
defparam \LessThan0~0 .lut_mask = 16'hFFFE;
defparam \LessThan0~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \LessThan0~1 (
	.dataa(b_full1),
	.datab(counter_reg_bit_5),
	.datac(counter_reg_bit_4),
	.datad(\LessThan0~0_combout ),
	.cin(gnd),
	.combout(\LessThan0~1_combout ),
	.cout());
defparam \LessThan0~1 .lut_mask = 16'h7FFF;
defparam \LessThan0~1 .sum_lutc_input = "datac";

dffeas fifo_AE(
	.clk(clk_clk),
	.d(\LessThan0~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_AE~q ),
	.prn(vcc));
defparam fifo_AE.is_wysiwyg = "true";
defparam fifo_AE.power_up = "low";

dffeas ien_AE(
	.clk(clk_clk),
	.d(src_payload2),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ien_AE~0_combout ),
	.q(\ien_AE~q ),
	.prn(vcc));
defparam ien_AE.is_wysiwyg = "true";
defparam ien_AE.power_up = "low";

cyclone10lp_lcell_comb \pause_irq~0 (
	.dataa(b_non_empty),
	.datab(\processor_jtag_uart_0_alt_jtag_atlantic|t_pause~reg0_q ),
	.datac(\pause_irq~q ),
	.datad(read_01),
	.cin(gnd),
	.combout(\pause_irq~0_combout ),
	.cout());
defparam \pause_irq~0 .lut_mask = 16'hFEFF;
defparam \pause_irq~0 .sum_lutc_input = "datac";

dffeas pause_irq(
	.clk(clk_clk),
	.d(\pause_irq~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pause_irq~q ),
	.prn(vcc));
defparam pause_irq.is_wysiwyg = "true";
defparam pause_irq.power_up = "low";

cyclone10lp_lcell_comb \Add0~0 (
	.dataa(counter_reg_bit_01),
	.datab(counter_reg_bit_11),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout(\Add0~1 ));
defparam \Add0~0 .lut_mask = 16'h6677;
defparam \Add0~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Add0~2 (
	.dataa(counter_reg_bit_21),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1 ),
	.combout(\Add0~2_combout ),
	.cout(\Add0~3 ));
defparam \Add0~2 .lut_mask = 16'h5AAF;
defparam \Add0~2 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add0~4 (
	.dataa(counter_reg_bit_31),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~3 ),
	.combout(\Add0~4_combout ),
	.cout(\Add0~5 ));
defparam \Add0~4 .lut_mask = 16'h5A5F;
defparam \Add0~4 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \LessThan1~0 (
	.dataa(\Add0~4_combout ),
	.datab(counter_reg_bit_01),
	.datac(\Add0~0_combout ),
	.datad(\Add0~2_combout ),
	.cin(gnd),
	.combout(\LessThan1~0_combout ),
	.cout());
defparam \LessThan1~0 .lut_mask = 16'hFFFE;
defparam \LessThan1~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Add0~6 (
	.dataa(counter_reg_bit_41),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~5 ),
	.combout(\Add0~6_combout ),
	.cout(\Add0~7 ));
defparam \Add0~6 .lut_mask = 16'h5AAF;
defparam \Add0~6 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add0~8 (
	.dataa(counter_reg_bit_51),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~7 ),
	.combout(\Add0~8_combout ),
	.cout(\Add0~9 ));
defparam \Add0~8 .lut_mask = 16'h5A5F;
defparam \Add0~8 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \LessThan1~1 (
	.dataa(\Add0~6_combout ),
	.datab(\Add0~8_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\LessThan1~1_combout ),
	.cout());
defparam \LessThan1~1 .lut_mask = 16'hEEEE;
defparam \LessThan1~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Add0~10 (
	.dataa(b_full),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~9 ),
	.combout(\Add0~10_combout ),
	.cout(\Add0~11 ));
defparam \Add0~10 .lut_mask = 16'h5AAF;
defparam \Add0~10 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add0~12 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add0~11 ),
	.combout(\Add0~12_combout ),
	.cout());
defparam \Add0~12 .lut_mask = 16'hF0F0;
defparam \Add0~12 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \LessThan1~2 (
	.dataa(\LessThan1~0_combout ),
	.datab(\LessThan1~1_combout ),
	.datac(\Add0~10_combout ),
	.datad(\Add0~12_combout ),
	.cin(gnd),
	.combout(\LessThan1~2_combout ),
	.cout());
defparam \LessThan1~2 .lut_mask = 16'h7FFF;
defparam \LessThan1~2 .sum_lutc_input = "datac";

dffeas fifo_AF(
	.clk(clk_clk),
	.d(\LessThan1~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_AF~q ),
	.prn(vcc));
defparam fifo_AF.is_wysiwyg = "true";
defparam fifo_AF.power_up = "low";

cyclone10lp_lcell_comb \woverflow~0 (
	.dataa(uav_write),
	.datab(saved_grant_0),
	.datac(\fifo_rd~0_combout ),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\woverflow~0_combout ),
	.cout());
defparam \woverflow~0 .lut_mask = 16'hFEFF;
defparam \woverflow~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \woverflow~1 (
	.dataa(b_full1),
	.datab(woverflow1),
	.datac(gnd),
	.datad(\woverflow~0_combout ),
	.cin(gnd),
	.combout(\woverflow~1_combout ),
	.cout());
defparam \woverflow~1 .lut_mask = 16'hAACC;
defparam \woverflow~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \rvalid~0 (
	.dataa(b_non_empty),
	.datab(rvalid1),
	.datac(gnd),
	.datad(\fifo_rd~2_combout ),
	.cin(gnd),
	.combout(\rvalid~0_combout ),
	.cout());
defparam \rvalid~0 .lut_mask = 16'hAACC;
defparam \rvalid~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ac~0 (
	.dataa(\processor_jtag_uart_0_alt_jtag_atlantic|t_ena~reg0_q ),
	.datab(\processor_jtag_uart_0_alt_jtag_atlantic|t_pause~reg0_q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ac~0_combout ),
	.cout());
defparam \ac~0 .lut_mask = 16'hEEEE;
defparam \ac~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ac~1 (
	.dataa(\ac~0_combout ),
	.datab(ac1),
	.datac(d_writedata_10),
	.datad(\ien_AE~0_combout ),
	.cin(gnd),
	.combout(\ac~1_combout ),
	.cout());
defparam \ac~1 .lut_mask = 16'hEFFF;
defparam \ac~1 .sum_lutc_input = "datac";

endmodule

module processor_alt_jtag_atlantic (
	r_dat,
	adapted_tdo1,
	rst_n,
	rst11,
	t_dav,
	rvalid01,
	r_val,
	r_ena11,
	t_ena,
	wdata_0,
	t_pause,
	wdata_1,
	wdata_4,
	wdata_3,
	wdata_2,
	wdata_5,
	wdata_7,
	wdata_6,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	splitter_nodes_receive_0_3,
	virtual_ir_scan_reg,
	clr_reg,
	state_3,
	state_8,
	irf_reg_0_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[7:0] r_dat;
output 	adapted_tdo1;
input 	rst_n;
output 	rst11;
input 	t_dav;
output 	rvalid01;
input 	r_val;
output 	r_ena11;
output 	t_ena;
output 	wdata_0;
output 	t_pause;
output 	wdata_1;
output 	wdata_4;
output 	wdata_3;
output 	wdata_2;
output 	wdata_5;
output 	wdata_7;
output 	wdata_6;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	splitter_nodes_receive_0_3;
input 	virtual_ir_scan_reg;
input 	clr_reg;
input 	state_3;
input 	state_8;
input 	irf_reg_0_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tck_t_dav~0_combout ;
wire \tck_t_dav~q ;
wire \state~1_combout ;
wire \always0~0_combout ;
wire \state~0_combout ;
wire \state~2_combout ;
wire \state~q ;
wire \count~9_combout ;
wire \td_shift[0]~4_combout ;
wire \count[2]~q ;
wire \count~8_combout ;
wire \count[3]~q ;
wire \count~7_combout ;
wire \count[4]~q ;
wire \count~6_combout ;
wire \count[5]~q ;
wire \count~5_combout ;
wire \count[6]~q ;
wire \count~4_combout ;
wire \count[7]~q ;
wire \count~2_combout ;
wire \count[8]~q ;
wire \count[9]~0_combout ;
wire \count[9]~q ;
wire \count~3_combout ;
wire \count[0]~q ;
wire \count~1_combout ;
wire \count[1]~q ;
wire \wdata[5]~2_combout ;
wire \user_saw_rvalid~0_combout ;
wire \user_saw_rvalid~q ;
wire \td_shift~10_combout ;
wire \td_shift[10]~q ;
wire \r_ena~0_combout ;
wire \rdata[7]~q ;
wire \td_shift~7_combout ;
wire \td_shift[9]~q ;
wire \td_shift~1_combout ;
wire \td_shift~11_combout ;
wire \rdata[6]~q ;
wire \td_shift~16_combout ;
wire \td_shift[8]~q ;
wire \rdata[5]~q ;
wire \td_shift~17_combout ;
wire \td_shift[7]~q ;
wire \rdata[4]~q ;
wire \td_shift~18_combout ;
wire \td_shift~19_combout ;
wire \td_shift[6]~q ;
wire \rdata[3]~q ;
wire \td_shift~14_combout ;
wire \td_shift~15_combout ;
wire \td_shift[5]~q ;
wire \rdata[2]~q ;
wire \td_shift~13_combout ;
wire \td_shift[4]~q ;
wire \rdata[1]~q ;
wire \td_shift~12_combout ;
wire \td_shift[3]~q ;
wire \rdata[0]~q ;
wire \td_shift~8_combout ;
wire \td_shift~9_combout ;
wire \td_shift[2]~q ;
wire \write_stalled~2_combout ;
wire \write_stalled~4_combout ;
wire \write_stalled~3_combout ;
wire \write_stalled~q ;
wire \td_shift~5_combout ;
wire \td_shift~6_combout ;
wire \td_shift[1]~q ;
wire \rvalid~q ;
wire \td_shift~0_combout ;
wire \td_shift~2_combout ;
wire \td_shift~3_combout ;
wire \td_shift[0]~q ;
wire \rvalid0~0_combout ;
wire \read~0_combout ;
wire \read~q ;
wire \read1~q ;
wire \read2~q ;
wire \read_req~q ;
wire \rvalid0~1_combout ;
wire \rst2~q ;
wire \rvalid0~2_combout ;
wire \write~0_combout ;
wire \wdata[5]~3_combout ;
wire \write~q ;
wire \write1~q ;
wire \write2~q ;
wire \write_valid~q ;
wire \t_ena~2_combout ;
wire \t_ena~3_combout ;
wire \always2~0_combout ;
wire \t_pause~0_combout ;
wire \jupdate~0_combout ;
wire \jupdate~q ;
wire \jupdate1~q ;
wire \jupdate2~q ;
wire \t_pause~1_combout ;


dffeas adapted_tdo(
	.clk(!altera_internal_jtag),
	.d(\td_shift[0]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(adapted_tdo1),
	.prn(vcc));
defparam adapted_tdo.is_wysiwyg = "true";
defparam adapted_tdo.power_up = "low";

dffeas rst1(
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rst11),
	.prn(vcc));
defparam rst1.is_wysiwyg = "true";
defparam rst1.power_up = "low";

dffeas rvalid0(
	.clk(clk),
	.d(\rvalid0~2_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rvalid01),
	.prn(vcc));
defparam rvalid0.is_wysiwyg = "true";
defparam rvalid0.power_up = "low";

dffeas r_ena1(
	.clk(clk),
	.d(\rvalid0~0_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_ena11),
	.prn(vcc));
defparam r_ena1.is_wysiwyg = "true";
defparam r_ena1.power_up = "low";

dffeas \t_ena~reg0 (
	.clk(clk),
	.d(\t_ena~3_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(t_ena),
	.prn(vcc));
defparam \t_ena~reg0 .is_wysiwyg = "true";
defparam \t_ena~reg0 .power_up = "low";

dffeas \wdata[0] (
	.clk(altera_internal_jtag),
	.d(altera_internal_jtag1),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~3_combout ),
	.q(wdata_0),
	.prn(vcc));
defparam \wdata[0] .is_wysiwyg = "true";
defparam \wdata[0] .power_up = "low";

dffeas \t_pause~reg0 (
	.clk(clk),
	.d(\t_pause~1_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(t_pause),
	.prn(vcc));
defparam \t_pause~reg0 .is_wysiwyg = "true";
defparam \t_pause~reg0 .power_up = "low";

dffeas \wdata[1] (
	.clk(altera_internal_jtag),
	.d(\td_shift[5]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[5]~3_combout ),
	.q(wdata_1),
	.prn(vcc));
defparam \wdata[1] .is_wysiwyg = "true";
defparam \wdata[1] .power_up = "low";

dffeas \wdata[4] (
	.clk(altera_internal_jtag),
	.d(\td_shift[8]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[5]~3_combout ),
	.q(wdata_4),
	.prn(vcc));
defparam \wdata[4] .is_wysiwyg = "true";
defparam \wdata[4] .power_up = "low";

dffeas \wdata[3] (
	.clk(altera_internal_jtag),
	.d(\td_shift[7]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[5]~3_combout ),
	.q(wdata_3),
	.prn(vcc));
defparam \wdata[3] .is_wysiwyg = "true";
defparam \wdata[3] .power_up = "low";

dffeas \wdata[2] (
	.clk(altera_internal_jtag),
	.d(\td_shift[6]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[5]~3_combout ),
	.q(wdata_2),
	.prn(vcc));
defparam \wdata[2] .is_wysiwyg = "true";
defparam \wdata[2] .power_up = "low";

dffeas \wdata[5] (
	.clk(altera_internal_jtag),
	.d(\td_shift[9]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[5]~3_combout ),
	.q(wdata_5),
	.prn(vcc));
defparam \wdata[5] .is_wysiwyg = "true";
defparam \wdata[5] .power_up = "low";

dffeas \wdata[7] (
	.clk(altera_internal_jtag),
	.d(altera_internal_jtag1),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[5]~3_combout ),
	.q(wdata_7),
	.prn(vcc));
defparam \wdata[7] .is_wysiwyg = "true";
defparam \wdata[7] .power_up = "low";

dffeas \wdata[6] (
	.clk(altera_internal_jtag),
	.d(\td_shift[10]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[5]~3_combout ),
	.q(wdata_6),
	.prn(vcc));
defparam \wdata[6] .is_wysiwyg = "true";
defparam \wdata[6] .power_up = "low";

cyclone10lp_lcell_comb \tck_t_dav~0 (
	.dataa(t_dav),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tck_t_dav~0_combout ),
	.cout());
defparam \tck_t_dav~0 .lut_mask = 16'h5555;
defparam \tck_t_dav~0 .sum_lutc_input = "datac";

dffeas tck_t_dav(
	.clk(altera_internal_jtag),
	.d(\tck_t_dav~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tck_t_dav~q ),
	.prn(vcc));
defparam tck_t_dav.is_wysiwyg = "true";
defparam tck_t_dav.power_up = "low";

cyclone10lp_lcell_comb \state~1 (
	.dataa(\state~q ),
	.datab(virtual_ir_scan_reg),
	.datac(splitter_nodes_receive_0_3),
	.datad(state_3),
	.cin(gnd),
	.combout(\state~1_combout ),
	.cout());
defparam \state~1 .lut_mask = 16'hEFFF;
defparam \state~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \always0~0 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(gnd),
	.datac(gnd),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
defparam \always0~0 .lut_mask = 16'hAAFF;
defparam \always0~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \state~0 (
	.dataa(altera_internal_jtag1),
	.datab(gnd),
	.datac(irf_reg_0_1),
	.datad(\state~q ),
	.cin(gnd),
	.combout(\state~0_combout ),
	.cout());
defparam \state~0 .lut_mask = 16'hAFFF;
defparam \state~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \state~2 (
	.dataa(\state~1_combout ),
	.datab(state_4),
	.datac(\always0~0_combout ),
	.datad(\state~0_combout ),
	.cin(gnd),
	.combout(\state~2_combout ),
	.cout());
defparam \state~2 .lut_mask = 16'hFFFE;
defparam \state~2 .sum_lutc_input = "datac";

dffeas state(
	.clk(altera_internal_jtag),
	.d(\state~2_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state~q ),
	.prn(vcc));
defparam state.is_wysiwyg = "true";
defparam state.power_up = "low";

cyclone10lp_lcell_comb \count~9 (
	.dataa(\count[1]~q ),
	.datab(state_4),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~9_combout ),
	.cout());
defparam \count~9 .lut_mask = 16'hEEEE;
defparam \count~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \td_shift[0]~4 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(state_4),
	.datac(state_3),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\td_shift[0]~4_combout ),
	.cout());
defparam \td_shift[0]~4 .lut_mask = 16'hFEFF;
defparam \td_shift[0]~4 .sum_lutc_input = "datac";

dffeas \count[2] (
	.clk(altera_internal_jtag),
	.d(\count~9_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[2]~q ),
	.prn(vcc));
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";

cyclone10lp_lcell_comb \count~8 (
	.dataa(state_4),
	.datab(\count[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~8_combout ),
	.cout());
defparam \count~8 .lut_mask = 16'hEEEE;
defparam \count~8 .sum_lutc_input = "datac";

dffeas \count[3] (
	.clk(altera_internal_jtag),
	.d(\count~8_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[3]~q ),
	.prn(vcc));
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";

cyclone10lp_lcell_comb \count~7 (
	.dataa(state_4),
	.datab(\count[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~7_combout ),
	.cout());
defparam \count~7 .lut_mask = 16'hEEEE;
defparam \count~7 .sum_lutc_input = "datac";

dffeas \count[4] (
	.clk(altera_internal_jtag),
	.d(\count~7_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[4]~q ),
	.prn(vcc));
defparam \count[4] .is_wysiwyg = "true";
defparam \count[4] .power_up = "low";

cyclone10lp_lcell_comb \count~6 (
	.dataa(state_4),
	.datab(\count[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~6_combout ),
	.cout());
defparam \count~6 .lut_mask = 16'hEEEE;
defparam \count~6 .sum_lutc_input = "datac";

dffeas \count[5] (
	.clk(altera_internal_jtag),
	.d(\count~6_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[5]~q ),
	.prn(vcc));
defparam \count[5] .is_wysiwyg = "true";
defparam \count[5] .power_up = "low";

cyclone10lp_lcell_comb \count~5 (
	.dataa(state_4),
	.datab(\count[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~5_combout ),
	.cout());
defparam \count~5 .lut_mask = 16'hEEEE;
defparam \count~5 .sum_lutc_input = "datac";

dffeas \count[6] (
	.clk(altera_internal_jtag),
	.d(\count~5_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[6]~q ),
	.prn(vcc));
defparam \count[6] .is_wysiwyg = "true";
defparam \count[6] .power_up = "low";

cyclone10lp_lcell_comb \count~4 (
	.dataa(state_4),
	.datab(\count[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~4_combout ),
	.cout());
defparam \count~4 .lut_mask = 16'hEEEE;
defparam \count~4 .sum_lutc_input = "datac";

dffeas \count[7] (
	.clk(altera_internal_jtag),
	.d(\count~4_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[7]~q ),
	.prn(vcc));
defparam \count[7] .is_wysiwyg = "true";
defparam \count[7] .power_up = "low";

cyclone10lp_lcell_comb \count~2 (
	.dataa(state_4),
	.datab(\count[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~2_combout ),
	.cout());
defparam \count~2 .lut_mask = 16'hEEEE;
defparam \count~2 .sum_lutc_input = "datac";

dffeas \count[8] (
	.clk(altera_internal_jtag),
	.d(\count~2_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[8]~q ),
	.prn(vcc));
defparam \count[8] .is_wysiwyg = "true";
defparam \count[8] .power_up = "low";

cyclone10lp_lcell_comb \count[9]~0 (
	.dataa(state_4),
	.datab(\state~0_combout ),
	.datac(\count[8]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\count[9]~0_combout ),
	.cout());
defparam \count[9]~0 .lut_mask = 16'h7F7F;
defparam \count[9]~0 .sum_lutc_input = "datac";

dffeas \count[9] (
	.clk(altera_internal_jtag),
	.d(\count[9]~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[9]~q ),
	.prn(vcc));
defparam \count[9] .is_wysiwyg = "true";
defparam \count[9] .power_up = "low";

cyclone10lp_lcell_comb \count~3 (
	.dataa(state_4),
	.datab(gnd),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\count~3_combout ),
	.cout());
defparam \count~3 .lut_mask = 16'hAAFF;
defparam \count~3 .sum_lutc_input = "datac";

dffeas \count[0] (
	.clk(altera_internal_jtag),
	.d(\count~3_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[0]~q ),
	.prn(vcc));
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";

cyclone10lp_lcell_comb \count~1 (
	.dataa(state_4),
	.datab(\count[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~1_combout ),
	.cout());
defparam \count~1 .lut_mask = 16'hEEEE;
defparam \count~1 .sum_lutc_input = "datac";

dffeas \count[1] (
	.clk(altera_internal_jtag),
	.d(\count~1_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[1]~q ),
	.prn(vcc));
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";

cyclone10lp_lcell_comb \wdata[5]~2 (
	.dataa(\state~q ),
	.datab(state_4),
	.datac(\always0~0_combout ),
	.datad(irf_reg_0_1),
	.cin(gnd),
	.combout(\wdata[5]~2_combout ),
	.cout());
defparam \wdata[5]~2 .lut_mask = 16'hFEFF;
defparam \wdata[5]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \user_saw_rvalid~0 (
	.dataa(\td_shift[0]~q ),
	.datab(\user_saw_rvalid~q ),
	.datac(\count[0]~q ),
	.datad(\wdata[5]~2_combout ),
	.cin(gnd),
	.combout(\user_saw_rvalid~0_combout ),
	.cout());
defparam \user_saw_rvalid~0 .lut_mask = 16'hEFFE;
defparam \user_saw_rvalid~0 .sum_lutc_input = "datac";

dffeas user_saw_rvalid(
	.clk(altera_internal_jtag),
	.d(\user_saw_rvalid~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\user_saw_rvalid~q ),
	.prn(vcc));
defparam user_saw_rvalid.is_wysiwyg = "true";
defparam user_saw_rvalid.power_up = "low";

cyclone10lp_lcell_comb \td_shift~10 (
	.dataa(altera_internal_jtag1),
	.datab(state_4),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\td_shift~10_combout ),
	.cout());
defparam \td_shift~10 .lut_mask = 16'hEEEE;
defparam \td_shift~10 .sum_lutc_input = "datac";

dffeas \td_shift[10] (
	.clk(altera_internal_jtag),
	.d(\td_shift~10_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[10]~q ),
	.prn(vcc));
defparam \td_shift[10] .is_wysiwyg = "true";
defparam \td_shift[10] .power_up = "low";

cyclone10lp_lcell_comb \r_ena~0 (
	.dataa(r_val),
	.datab(r_ena11),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\r_ena~0_combout ),
	.cout());
defparam \r_ena~0 .lut_mask = 16'hEEEE;
defparam \r_ena~0 .sum_lutc_input = "datac";

dffeas \rdata[7] (
	.clk(clk),
	.d(r_dat[7]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[7]~q ),
	.prn(vcc));
defparam \rdata[7] .is_wysiwyg = "true";
defparam \rdata[7] .power_up = "low";

cyclone10lp_lcell_comb \td_shift~7 (
	.dataa(\td_shift[10]~q ),
	.datab(\rdata[7]~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~7_combout ),
	.cout());
defparam \td_shift~7 .lut_mask = 16'hAACC;
defparam \td_shift~7 .sum_lutc_input = "datac";

dffeas \td_shift[9] (
	.clk(altera_internal_jtag),
	.d(\td_shift~7_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[9]~q ),
	.prn(vcc));
defparam \td_shift[9] .is_wysiwyg = "true";
defparam \td_shift[9] .power_up = "low";

cyclone10lp_lcell_comb \td_shift~1 (
	.dataa(\state~q ),
	.datab(\count[1]~q ),
	.datac(\user_saw_rvalid~q ),
	.datad(\td_shift[9]~q ),
	.cin(gnd),
	.combout(\td_shift~1_combout ),
	.cout());
defparam \td_shift~1 .lut_mask = 16'hEFFF;
defparam \td_shift~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \td_shift~11 (
	.dataa(state_4),
	.datab(irf_reg_0_1),
	.datac(gnd),
	.datad(\td_shift~1_combout ),
	.cin(gnd),
	.combout(\td_shift~11_combout ),
	.cout());
defparam \td_shift~11 .lut_mask = 16'hEEFF;
defparam \td_shift~11 .sum_lutc_input = "datac";

dffeas \rdata[6] (
	.clk(clk),
	.d(r_dat[6]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[6]~q ),
	.prn(vcc));
defparam \rdata[6] .is_wysiwyg = "true";
defparam \rdata[6] .power_up = "low";

cyclone10lp_lcell_comb \td_shift~16 (
	.dataa(\td_shift[9]~q ),
	.datab(\rdata[6]~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~16_combout ),
	.cout());
defparam \td_shift~16 .lut_mask = 16'hAACC;
defparam \td_shift~16 .sum_lutc_input = "datac";

dffeas \td_shift[8] (
	.clk(altera_internal_jtag),
	.d(\td_shift~16_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[8]~q ),
	.prn(vcc));
defparam \td_shift[8] .is_wysiwyg = "true";
defparam \td_shift[8] .power_up = "low";

dffeas \rdata[5] (
	.clk(clk),
	.d(r_dat[5]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[5]~q ),
	.prn(vcc));
defparam \rdata[5] .is_wysiwyg = "true";
defparam \rdata[5] .power_up = "low";

cyclone10lp_lcell_comb \td_shift~17 (
	.dataa(\td_shift~11_combout ),
	.datab(\td_shift[8]~q ),
	.datac(\rdata[5]~q ),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~17_combout ),
	.cout());
defparam \td_shift~17 .lut_mask = 16'hFAFC;
defparam \td_shift~17 .sum_lutc_input = "datac";

dffeas \td_shift[7] (
	.clk(altera_internal_jtag),
	.d(\td_shift~17_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[7]~q ),
	.prn(vcc));
defparam \td_shift[7] .is_wysiwyg = "true";
defparam \td_shift[7] .power_up = "low";

dffeas \rdata[4] (
	.clk(clk),
	.d(r_dat[4]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[4]~q ),
	.prn(vcc));
defparam \rdata[4] .is_wysiwyg = "true";
defparam \rdata[4] .power_up = "low";

cyclone10lp_lcell_comb \td_shift~18 (
	.dataa(\td_shift[7]~q ),
	.datab(\rdata[4]~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~18_combout ),
	.cout());
defparam \td_shift~18 .lut_mask = 16'hAACC;
defparam \td_shift~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \td_shift~19 (
	.dataa(irf_reg_0_1),
	.datab(\td_shift~18_combout ),
	.datac(state_4),
	.datad(\td_shift~1_combout ),
	.cin(gnd),
	.combout(\td_shift~19_combout ),
	.cout());
defparam \td_shift~19 .lut_mask = 16'hACFF;
defparam \td_shift~19 .sum_lutc_input = "datac";

dffeas \td_shift[6] (
	.clk(altera_internal_jtag),
	.d(\td_shift~19_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[6]~q ),
	.prn(vcc));
defparam \td_shift[6] .is_wysiwyg = "true";
defparam \td_shift[6] .power_up = "low";

dffeas \rdata[3] (
	.clk(clk),
	.d(r_dat[3]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[3]~q ),
	.prn(vcc));
defparam \rdata[3] .is_wysiwyg = "true";
defparam \rdata[3] .power_up = "low";

cyclone10lp_lcell_comb \td_shift~14 (
	.dataa(\td_shift[6]~q ),
	.datab(\rdata[3]~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~14_combout ),
	.cout());
defparam \td_shift~14 .lut_mask = 16'hAACC;
defparam \td_shift~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \td_shift~15 (
	.dataa(irf_reg_0_1),
	.datab(\td_shift~14_combout ),
	.datac(state_4),
	.datad(\td_shift~1_combout ),
	.cin(gnd),
	.combout(\td_shift~15_combout ),
	.cout());
defparam \td_shift~15 .lut_mask = 16'hACFF;
defparam \td_shift~15 .sum_lutc_input = "datac";

dffeas \td_shift[5] (
	.clk(altera_internal_jtag),
	.d(\td_shift~15_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[5]~q ),
	.prn(vcc));
defparam \td_shift[5] .is_wysiwyg = "true";
defparam \td_shift[5] .power_up = "low";

dffeas \rdata[2] (
	.clk(clk),
	.d(r_dat[2]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[2]~q ),
	.prn(vcc));
defparam \rdata[2] .is_wysiwyg = "true";
defparam \rdata[2] .power_up = "low";

cyclone10lp_lcell_comb \td_shift~13 (
	.dataa(\td_shift~11_combout ),
	.datab(\td_shift[5]~q ),
	.datac(\rdata[2]~q ),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~13_combout ),
	.cout());
defparam \td_shift~13 .lut_mask = 16'hFAFC;
defparam \td_shift~13 .sum_lutc_input = "datac";

dffeas \td_shift[4] (
	.clk(altera_internal_jtag),
	.d(\td_shift~13_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[4]~q ),
	.prn(vcc));
defparam \td_shift[4] .is_wysiwyg = "true";
defparam \td_shift[4] .power_up = "low";

dffeas \rdata[1] (
	.clk(clk),
	.d(r_dat[1]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[1]~q ),
	.prn(vcc));
defparam \rdata[1] .is_wysiwyg = "true";
defparam \rdata[1] .power_up = "low";

cyclone10lp_lcell_comb \td_shift~12 (
	.dataa(\td_shift~11_combout ),
	.datab(\td_shift[4]~q ),
	.datac(\rdata[1]~q ),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~12_combout ),
	.cout());
defparam \td_shift~12 .lut_mask = 16'hFAFC;
defparam \td_shift~12 .sum_lutc_input = "datac";

dffeas \td_shift[3] (
	.clk(altera_internal_jtag),
	.d(\td_shift~12_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[3]~q ),
	.prn(vcc));
defparam \td_shift[3] .is_wysiwyg = "true";
defparam \td_shift[3] .power_up = "low";

dffeas \rdata[0] (
	.clk(clk),
	.d(r_dat[0]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[0]~q ),
	.prn(vcc));
defparam \rdata[0] .is_wysiwyg = "true";
defparam \rdata[0] .power_up = "low";

cyclone10lp_lcell_comb \td_shift~8 (
	.dataa(\td_shift[3]~q ),
	.datab(\rdata[0]~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~8_combout ),
	.cout());
defparam \td_shift~8 .lut_mask = 16'hAACC;
defparam \td_shift~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \td_shift~9 (
	.dataa(irf_reg_0_1),
	.datab(\td_shift~8_combout ),
	.datac(state_4),
	.datad(\td_shift~1_combout ),
	.cin(gnd),
	.combout(\td_shift~9_combout ),
	.cout());
defparam \td_shift~9 .lut_mask = 16'hACFF;
defparam \td_shift~9 .sum_lutc_input = "datac";

dffeas \td_shift[2] (
	.clk(altera_internal_jtag),
	.d(\td_shift~9_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[2]~q ),
	.prn(vcc));
defparam \td_shift[2] .is_wysiwyg = "true";
defparam \td_shift[2] .power_up = "low";

cyclone10lp_lcell_comb \write_stalled~2 (
	.dataa(\write_stalled~q ),
	.datab(\td_shift[10]~q ),
	.datac(altera_internal_jtag1),
	.datad(\tck_t_dav~q ),
	.cin(gnd),
	.combout(\write_stalled~2_combout ),
	.cout());
defparam \write_stalled~2 .lut_mask = 16'hEFFF;
defparam \write_stalled~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \write_stalled~4 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(virtual_ir_scan_reg),
	.datac(irf_reg_0_1),
	.datad(gnd),
	.cin(gnd),
	.combout(\write_stalled~4_combout ),
	.cout());
defparam \write_stalled~4 .lut_mask = 16'hBFBF;
defparam \write_stalled~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \write_stalled~3 (
	.dataa(\count[1]~q ),
	.datab(\state~q ),
	.datac(state_4),
	.datad(\write_stalled~4_combout ),
	.cin(gnd),
	.combout(\write_stalled~3_combout ),
	.cout());
defparam \write_stalled~3 .lut_mask = 16'hFFFE;
defparam \write_stalled~3 .sum_lutc_input = "datac";

dffeas write_stalled(
	.clk(altera_internal_jtag),
	.d(\write_stalled~2_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~3_combout ),
	.q(\write_stalled~q ),
	.prn(vcc));
defparam write_stalled.is_wysiwyg = "true";
defparam write_stalled.power_up = "low";

cyclone10lp_lcell_comb \td_shift~5 (
	.dataa(\td_shift[2]~q ),
	.datab(\write_stalled~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~5_combout ),
	.cout());
defparam \td_shift~5 .lut_mask = 16'hAACC;
defparam \td_shift~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \td_shift~6 (
	.dataa(irf_reg_0_1),
	.datab(\td_shift~5_combout ),
	.datac(state_4),
	.datad(\td_shift~1_combout ),
	.cin(gnd),
	.combout(\td_shift~6_combout ),
	.cout());
defparam \td_shift~6 .lut_mask = 16'hACFF;
defparam \td_shift~6 .sum_lutc_input = "datac";

dffeas \td_shift[1] (
	.clk(altera_internal_jtag),
	.d(\td_shift~6_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[1]~q ),
	.prn(vcc));
defparam \td_shift[1] .is_wysiwyg = "true";
defparam \td_shift[1] .power_up = "low";

dffeas rvalid(
	.clk(clk),
	.d(rvalid01),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rvalid~q ),
	.prn(vcc));
defparam rvalid.is_wysiwyg = "true";
defparam rvalid.power_up = "low";

cyclone10lp_lcell_comb \td_shift~0 (
	.dataa(\td_shift[1]~q ),
	.datab(\rvalid~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~0_combout ),
	.cout());
defparam \td_shift~0 .lut_mask = 16'hAACC;
defparam \td_shift~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \td_shift~2 (
	.dataa(\td_shift~1_combout ),
	.datab(altera_internal_jtag1),
	.datac(\state~q ),
	.datad(irf_reg_0_1),
	.cin(gnd),
	.combout(\td_shift~2_combout ),
	.cout());
defparam \td_shift~2 .lut_mask = 16'hEFFF;
defparam \td_shift~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \td_shift~3 (
	.dataa(\tck_t_dav~q ),
	.datab(\td_shift~0_combout ),
	.datac(\td_shift~2_combout ),
	.datad(\state~q ),
	.cin(gnd),
	.combout(\td_shift~3_combout ),
	.cout());
defparam \td_shift~3 .lut_mask = 16'hACFF;
defparam \td_shift~3 .sum_lutc_input = "datac";

dffeas \td_shift[0] (
	.clk(altera_internal_jtag),
	.d(\td_shift~3_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[0]~q ),
	.prn(vcc));
defparam \td_shift[0] .is_wysiwyg = "true";
defparam \td_shift[0] .power_up = "low";

cyclone10lp_lcell_comb \rvalid0~0 (
	.dataa(rvalid01),
	.datab(r_val),
	.datac(r_ena11),
	.datad(gnd),
	.cin(gnd),
	.combout(\rvalid0~0_combout ),
	.cout());
defparam \rvalid0~0 .lut_mask = 16'h7F7F;
defparam \rvalid0~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \read~0 (
	.dataa(\read~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\read~0_combout ),
	.cout());
defparam \read~0 .lut_mask = 16'h5555;
defparam \read~0 .sum_lutc_input = "datac";

dffeas read(
	.clk(altera_internal_jtag),
	.d(\read~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~3_combout ),
	.q(\read~q ),
	.prn(vcc));
defparam read.is_wysiwyg = "true";
defparam read.power_up = "low";

dffeas read1(
	.clk(clk),
	.d(\read~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read1~q ),
	.prn(vcc));
defparam read1.is_wysiwyg = "true";
defparam read1.power_up = "low";

dffeas read2(
	.clk(clk),
	.d(\read1~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read2~q ),
	.prn(vcc));
defparam read2.is_wysiwyg = "true";
defparam read2.power_up = "low";

dffeas read_req(
	.clk(altera_internal_jtag),
	.d(\td_shift[9]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~3_combout ),
	.q(\read_req~q ),
	.prn(vcc));
defparam read_req.is_wysiwyg = "true";
defparam read_req.power_up = "low";

cyclone10lp_lcell_comb \rvalid0~1 (
	.dataa(\read1~q ),
	.datab(\read2~q ),
	.datac(\user_saw_rvalid~q ),
	.datad(\read_req~q ),
	.cin(gnd),
	.combout(\rvalid0~1_combout ),
	.cout());
defparam \rvalid0~1 .lut_mask = 16'h6FFF;
defparam \rvalid0~1 .sum_lutc_input = "datac";

dffeas rst2(
	.clk(clk),
	.d(rst11),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rst2~q ),
	.prn(vcc));
defparam rst2.is_wysiwyg = "true";
defparam rst2.power_up = "low";

cyclone10lp_lcell_comb \rvalid0~2 (
	.dataa(\rvalid0~0_combout ),
	.datab(\rvalid0~1_combout ),
	.datac(gnd),
	.datad(\rst2~q ),
	.cin(gnd),
	.combout(\rvalid0~2_combout ),
	.cout());
defparam \rvalid0~2 .lut_mask = 16'hDDFF;
defparam \rvalid0~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \write~0 (
	.dataa(\write~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\write~0_combout ),
	.cout());
defparam \write~0 .lut_mask = 16'h5555;
defparam \write~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wdata[5]~3 (
	.dataa(\count[8]~q ),
	.datab(\state~q ),
	.datac(state_4),
	.datad(\write_stalled~4_combout ),
	.cin(gnd),
	.combout(\wdata[5]~3_combout ),
	.cout());
defparam \wdata[5]~3 .lut_mask = 16'hFFFE;
defparam \wdata[5]~3 .sum_lutc_input = "datac";

dffeas write(
	.clk(altera_internal_jtag),
	.d(\write~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[5]~3_combout ),
	.q(\write~q ),
	.prn(vcc));
defparam write.is_wysiwyg = "true";
defparam write.power_up = "low";

dffeas write1(
	.clk(clk),
	.d(\write~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write1~q ),
	.prn(vcc));
defparam write1.is_wysiwyg = "true";
defparam write1.power_up = "low";

dffeas write2(
	.clk(clk),
	.d(\write1~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write2~q ),
	.prn(vcc));
defparam write2.is_wysiwyg = "true";
defparam write2.power_up = "low";

dffeas write_valid(
	.clk(altera_internal_jtag),
	.d(\td_shift[10]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~3_combout ),
	.q(\write_valid~q ),
	.prn(vcc));
defparam write_valid.is_wysiwyg = "true";
defparam write_valid.power_up = "low";

cyclone10lp_lcell_comb \t_ena~2 (
	.dataa(t_ena),
	.datab(\write_valid~q ),
	.datac(t_dav),
	.datad(\write_stalled~q ),
	.cin(gnd),
	.combout(\t_ena~2_combout ),
	.cout());
defparam \t_ena~2 .lut_mask = 16'hEFFF;
defparam \t_ena~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \t_ena~3 (
	.dataa(\write1~q ),
	.datab(\write2~q ),
	.datac(\rst2~q ),
	.datad(\t_ena~2_combout ),
	.cin(gnd),
	.combout(\t_ena~3_combout ),
	.cout());
defparam \t_ena~3 .lut_mask = 16'hFFF6;
defparam \t_ena~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \always2~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\write1~q ),
	.datad(\write2~q ),
	.cin(gnd),
	.combout(\always2~0_combout ),
	.cout());
defparam \always2~0 .lut_mask = 16'h0FF0;
defparam \always2~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \t_pause~0 (
	.dataa(\always2~0_combout ),
	.datab(t_dav),
	.datac(\write_stalled~q ),
	.datad(\write_valid~q ),
	.cin(gnd),
	.combout(\t_pause~0_combout ),
	.cout());
defparam \t_pause~0 .lut_mask = 16'hFEFF;
defparam \t_pause~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \jupdate~0 (
	.dataa(\jupdate~q ),
	.datab(irf_reg_0_1),
	.datac(\always0~0_combout ),
	.datad(state_8),
	.cin(gnd),
	.combout(\jupdate~0_combout ),
	.cout());
defparam \jupdate~0 .lut_mask = 16'h6996;
defparam \jupdate~0 .sum_lutc_input = "datac";

dffeas jupdate(
	.clk(!altera_internal_jtag),
	.d(\jupdate~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jupdate~q ),
	.prn(vcc));
defparam jupdate.is_wysiwyg = "true";
defparam jupdate.power_up = "low";

dffeas jupdate1(
	.clk(clk),
	.d(\jupdate~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jupdate1~q ),
	.prn(vcc));
defparam jupdate1.is_wysiwyg = "true";
defparam jupdate1.power_up = "low";

dffeas jupdate2(
	.clk(clk),
	.d(\jupdate1~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jupdate2~q ),
	.prn(vcc));
defparam jupdate2.is_wysiwyg = "true";
defparam jupdate2.power_up = "low";

cyclone10lp_lcell_comb \t_pause~1 (
	.dataa(\rst2~q ),
	.datab(\t_pause~0_combout ),
	.datac(\jupdate1~q ),
	.datad(\jupdate2~q ),
	.cin(gnd),
	.combout(\t_pause~1_combout ),
	.cout());
defparam \t_pause~1 .lut_mask = 16'hEFFE;
defparam \t_pause~1 .sum_lutc_input = "datac";

endmodule

module processor_processor_jtag_uart_0_scfifo_r (
	q_b_0,
	q_b_1,
	q_b_4,
	q_b_3,
	q_b_2,
	q_b_5,
	q_b_7,
	q_b_6,
	r_sync_rst,
	b_full,
	counter_reg_bit_0,
	b_non_empty,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	t_ena,
	fifo_rd,
	wr_rfifo,
	wdata_0,
	fifo_rd1,
	wdata_1,
	wdata_4,
	wdata_3,
	wdata_2,
	wdata_5,
	wdata_7,
	wdata_6,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_0;
output 	q_b_1;
output 	q_b_4;
output 	q_b_3;
output 	q_b_2;
output 	q_b_5;
output 	q_b_7;
output 	q_b_6;
input 	r_sync_rst;
output 	b_full;
output 	counter_reg_bit_0;
output 	b_non_empty;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
input 	t_ena;
input 	fifo_rd;
input 	wr_rfifo;
input 	wdata_0;
input 	fifo_rd1;
input 	wdata_1;
input 	wdata_4;
input 	wdata_3;
input 	wdata_2;
input 	wdata_5;
input 	wdata_7;
input 	wdata_6;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



processor_scfifo_1 rfifo(
	.q({q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.r_sync_rst(r_sync_rst),
	.b_full(b_full),
	.counter_reg_bit_0(counter_reg_bit_0),
	.b_non_empty(b_non_empty),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.t_ena(t_ena),
	.fifo_rd(fifo_rd),
	.wrreq(wr_rfifo),
	.data({wdata_7,wdata_6,wdata_5,wdata_4,wdata_3,wdata_2,wdata_1,wdata_0}),
	.fifo_rd1(fifo_rd1),
	.clock(clk_clk));

endmodule

module processor_scfifo_1 (
	q,
	r_sync_rst,
	b_full,
	counter_reg_bit_0,
	b_non_empty,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	t_ena,
	fifo_rd,
	wrreq,
	data,
	fifo_rd1,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	r_sync_rst;
output 	b_full;
output 	counter_reg_bit_0;
output 	b_non_empty;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
input 	t_ena;
input 	fifo_rd;
input 	wrreq;
input 	[7:0] data;
input 	fifo_rd1;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



processor_scfifo_cr21 auto_generated(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.r_sync_rst(r_sync_rst),
	.b_full(b_full),
	.counter_reg_bit_0(counter_reg_bit_0),
	.b_non_empty(b_non_empty),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.t_ena(t_ena),
	.fifo_rd(fifo_rd),
	.wrreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.fifo_rd1(fifo_rd1),
	.clock(clock));

endmodule

module processor_scfifo_cr21 (
	q,
	r_sync_rst,
	b_full,
	counter_reg_bit_0,
	b_non_empty,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	t_ena,
	fifo_rd,
	wrreq,
	data,
	fifo_rd1,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	r_sync_rst;
output 	b_full;
output 	counter_reg_bit_0;
output 	b_non_empty;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
input 	t_ena;
input 	fifo_rd;
input 	wrreq;
input 	[7:0] data;
input 	fifo_rd1;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



processor_a_dpfifo_e011 dpfifo(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.r_sync_rst(r_sync_rst),
	.b_full(b_full),
	.counter_reg_bit_0(counter_reg_bit_0),
	.b_non_empty(b_non_empty),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.t_ena(t_ena),
	.fifo_rd(fifo_rd),
	.wreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.fifo_rd1(fifo_rd1),
	.clock(clock));

endmodule

module processor_a_dpfifo_e011 (
	q,
	r_sync_rst,
	b_full,
	counter_reg_bit_0,
	b_non_empty,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	t_ena,
	fifo_rd,
	wreq,
	data,
	fifo_rd1,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	r_sync_rst;
output 	b_full;
output 	counter_reg_bit_0;
output 	b_non_empty;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
input 	t_ena;
input 	fifo_rd;
input 	wreq;
input 	[7:0] data;
input 	fifo_rd1;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \wr_ptr|counter_reg_bit[5]~q ;
wire \rd_ptr_count|counter_reg_bit[0]~q ;
wire \rd_ptr_count|counter_reg_bit[1]~q ;
wire \rd_ptr_count|counter_reg_bit[2]~q ;
wire \rd_ptr_count|counter_reg_bit[3]~q ;
wire \rd_ptr_count|counter_reg_bit[4]~q ;
wire \rd_ptr_count|counter_reg_bit[5]~q ;


processor_cntr_qnb_1 wr_ptr(
	.r_sync_rst(r_sync_rst),
	.wr_rfifo(wreq),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\wr_ptr|counter_reg_bit[5]~q ),
	.clock(clock));

processor_cntr_qnb rd_ptr_count(
	.r_sync_rst(r_sync_rst),
	.fifo_rd(fifo_rd),
	.counter_reg_bit_0(\rd_ptr_count|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_count|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_count|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_count|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\rd_ptr_count|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\rd_ptr_count|counter_reg_bit[5]~q ),
	.clock(clock));

processor_altsyncram_gio1 FIFOram(
	.q_b({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.clocken1(fifo_rd),
	.wren_a(wreq),
	.data_a({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_a({\wr_ptr|counter_reg_bit[5]~q ,\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.address_b({\rd_ptr_count|counter_reg_bit[5]~q ,\rd_ptr_count|counter_reg_bit[4]~q ,\rd_ptr_count|counter_reg_bit[3]~q ,\rd_ptr_count|counter_reg_bit[2]~q ,\rd_ptr_count|counter_reg_bit[1]~q ,\rd_ptr_count|counter_reg_bit[0]~q }),
	.clock1(clock),
	.clock0(clock));

processor_a_fefifo_7cf fifo_state(
	.r_sync_rst(r_sync_rst),
	.b_full1(b_full),
	.counter_reg_bit_0(counter_reg_bit_0),
	.b_non_empty1(b_non_empty),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.t_ena(t_ena),
	.fifo_rd(fifo_rd),
	.wreq(wreq),
	.fifo_rd1(fifo_rd1),
	.clock(clock));

endmodule

module processor_a_fefifo_7cf (
	r_sync_rst,
	b_full1,
	counter_reg_bit_0,
	b_non_empty1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	t_ena,
	fifo_rd,
	wreq,
	fifo_rd1,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	b_full1;
output 	counter_reg_bit_0;
output 	b_non_empty1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
input 	t_ena;
input 	fifo_rd;
input 	wreq;
input 	fifo_rd1;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \_~4_combout ;
wire \b_full~0_combout ;
wire \b_full~1_combout ;
wire \b_full~2_combout ;
wire \b_non_empty~0_combout ;
wire \_~2_combout ;
wire \_~3_combout ;
wire \b_non_empty~1_combout ;


processor_cntr_6o7 count_usedw(
	.r_sync_rst(r_sync_rst),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.updown(wreq),
	._(\_~4_combout ),
	.clock(clock));

cyclone10lp_lcell_comb \_~4 (
	.dataa(t_ena),
	.datab(b_full1),
	.datac(b_non_empty1),
	.datad(fifo_rd1),
	.cin(gnd),
	.combout(\_~4_combout ),
	.cout());
defparam \_~4 .lut_mask = 16'h6996;
defparam \_~4 .sum_lutc_input = "datac";

dffeas b_full(
	.clk(clock),
	.d(\b_full~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_full1),
	.prn(vcc));
defparam b_full.is_wysiwyg = "true";
defparam b_full.power_up = "low";

dffeas b_non_empty(
	.clk(clock),
	.d(\b_non_empty~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_non_empty1),
	.prn(vcc));
defparam b_non_empty.is_wysiwyg = "true";
defparam b_non_empty.power_up = "low";

cyclone10lp_lcell_comb \b_full~0 (
	.dataa(b_non_empty1),
	.datab(counter_reg_bit_5),
	.datac(counter_reg_bit_4),
	.datad(counter_reg_bit_3),
	.cin(gnd),
	.combout(\b_full~0_combout ),
	.cout());
defparam \b_full~0 .lut_mask = 16'hFFFE;
defparam \b_full~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \b_full~1 (
	.dataa(counter_reg_bit_0),
	.datab(counter_reg_bit_2),
	.datac(counter_reg_bit_1),
	.datad(t_ena),
	.cin(gnd),
	.combout(\b_full~1_combout ),
	.cout());
defparam \b_full~1 .lut_mask = 16'hFFFE;
defparam \b_full~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \b_full~2 (
	.dataa(b_full1),
	.datab(\b_full~0_combout ),
	.datac(\b_full~1_combout ),
	.datad(fifo_rd),
	.cin(gnd),
	.combout(\b_full~2_combout ),
	.cout());
defparam \b_full~2 .lut_mask = 16'hFEFF;
defparam \b_full~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \b_non_empty~0 (
	.dataa(b_full1),
	.datab(t_ena),
	.datac(gnd),
	.datad(b_non_empty1),
	.cin(gnd),
	.combout(\b_non_empty~0_combout ),
	.cout());
defparam \b_non_empty~0 .lut_mask = 16'hEEFF;
defparam \b_non_empty~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_~2 (
	.dataa(counter_reg_bit_3),
	.datab(counter_reg_bit_2),
	.datac(counter_reg_bit_1),
	.datad(counter_reg_bit_0),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFEFF;
defparam \_~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_~3 (
	.dataa(counter_reg_bit_5),
	.datab(counter_reg_bit_4),
	.datac(wreq),
	.datad(\_~2_combout ),
	.cin(gnd),
	.combout(\_~3_combout ),
	.cout());
defparam \_~3 .lut_mask = 16'hFFFE;
defparam \_~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \b_non_empty~1 (
	.dataa(\b_non_empty~0_combout ),
	.datab(b_non_empty1),
	.datac(\_~3_combout ),
	.datad(fifo_rd1),
	.cin(gnd),
	.combout(\b_non_empty~1_combout ),
	.cout());
defparam \b_non_empty~1 .lut_mask = 16'hFEFF;
defparam \b_non_empty~1 .sum_lutc_input = "datac";

endmodule

module processor_cntr_6o7 (
	r_sync_rst,
	counter_reg_bit_0,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	updown,
	_,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	counter_reg_bit_0;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
input 	updown;
input 	_;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita1~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

cyclone10lp_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cyclone10lp_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cyclone10lp_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cyclone10lp_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cyclone10lp_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5A6F;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cyclone10lp_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module processor_altsyncram_gio1 (
	q_b,
	clocken1,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_b;
input 	clocken1;
input 	wren_a;
input 	[7:0] data_a;
input 	[5:0] address_a;
input 	[5:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

cyclone10lp_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk1_core_clock_enable = "ena1";
defparam ram_block1a0.clk1_input_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "processor_jtag_uart_0:jtag_uart_0|processor_jtag_uart_0_scfifo_r:the_processor_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_cr21:auto_generated|a_dpfifo_e011:dpfifo|altsyncram_gio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 6;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 63;
defparam ram_block1a0.port_a_logical_ram_depth = 64;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 6;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 63;
defparam ram_block1a0.port_b_logical_ram_depth = 64;
defparam ram_block1a0.port_b_logical_ram_width = 8;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk1_core_clock_enable = "ena1";
defparam ram_block1a1.clk1_input_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "processor_jtag_uart_0:jtag_uart_0|processor_jtag_uart_0_scfifo_r:the_processor_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_cr21:auto_generated|a_dpfifo_e011:dpfifo|altsyncram_gio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 6;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 63;
defparam ram_block1a1.port_a_logical_ram_depth = 64;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 6;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 63;
defparam ram_block1a1.port_b_logical_ram_depth = 64;
defparam ram_block1a1.port_b_logical_ram_width = 8;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk1_core_clock_enable = "ena1";
defparam ram_block1a4.clk1_input_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "processor_jtag_uart_0:jtag_uart_0|processor_jtag_uart_0_scfifo_r:the_processor_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_cr21:auto_generated|a_dpfifo_e011:dpfifo|altsyncram_gio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 6;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 63;
defparam ram_block1a4.port_a_logical_ram_depth = 64;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 6;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 63;
defparam ram_block1a4.port_b_logical_ram_depth = 64;
defparam ram_block1a4.port_b_logical_ram_width = 8;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk1_core_clock_enable = "ena1";
defparam ram_block1a3.clk1_input_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "processor_jtag_uart_0:jtag_uart_0|processor_jtag_uart_0_scfifo_r:the_processor_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_cr21:auto_generated|a_dpfifo_e011:dpfifo|altsyncram_gio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 6;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 63;
defparam ram_block1a3.port_a_logical_ram_depth = 64;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 6;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 63;
defparam ram_block1a3.port_b_logical_ram_depth = 64;
defparam ram_block1a3.port_b_logical_ram_width = 8;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk1_core_clock_enable = "ena1";
defparam ram_block1a2.clk1_input_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "processor_jtag_uart_0:jtag_uart_0|processor_jtag_uart_0_scfifo_r:the_processor_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_cr21:auto_generated|a_dpfifo_e011:dpfifo|altsyncram_gio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 6;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 63;
defparam ram_block1a2.port_a_logical_ram_depth = 64;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 6;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 63;
defparam ram_block1a2.port_b_logical_ram_depth = 64;
defparam ram_block1a2.port_b_logical_ram_width = 8;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk1_core_clock_enable = "ena1";
defparam ram_block1a5.clk1_input_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "processor_jtag_uart_0:jtag_uart_0|processor_jtag_uart_0_scfifo_r:the_processor_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_cr21:auto_generated|a_dpfifo_e011:dpfifo|altsyncram_gio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 6;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 63;
defparam ram_block1a5.port_a_logical_ram_depth = 64;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 6;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 63;
defparam ram_block1a5.port_b_logical_ram_depth = 64;
defparam ram_block1a5.port_b_logical_ram_width = 8;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk1_core_clock_enable = "ena1";
defparam ram_block1a7.clk1_input_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "processor_jtag_uart_0:jtag_uart_0|processor_jtag_uart_0_scfifo_r:the_processor_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_cr21:auto_generated|a_dpfifo_e011:dpfifo|altsyncram_gio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 6;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 63;
defparam ram_block1a7.port_a_logical_ram_depth = 64;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 6;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 63;
defparam ram_block1a7.port_b_logical_ram_depth = 64;
defparam ram_block1a7.port_b_logical_ram_width = 8;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk1_core_clock_enable = "ena1";
defparam ram_block1a6.clk1_input_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "processor_jtag_uart_0:jtag_uart_0|processor_jtag_uart_0_scfifo_r:the_processor_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_cr21:auto_generated|a_dpfifo_e011:dpfifo|altsyncram_gio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 6;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 63;
defparam ram_block1a6.port_a_logical_ram_depth = 64;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 6;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 63;
defparam ram_block1a6.port_b_logical_ram_depth = 64;
defparam ram_block1a6.port_b_logical_ram_width = 8;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

endmodule

module processor_cntr_qnb (
	r_sync_rst,
	fifo_rd,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	fifo_rd;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cyclone10lp_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cyclone10lp_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cyclone10lp_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cyclone10lp_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cyclone10lp_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cyclone10lp_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module processor_cntr_qnb_1 (
	r_sync_rst,
	wr_rfifo,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	wr_rfifo;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cyclone10lp_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cyclone10lp_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cyclone10lp_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cyclone10lp_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cyclone10lp_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cyclone10lp_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module processor_processor_jtag_uart_0_scfifo_w (
	q_b_7,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_6,
	q_b_5,
	q_b_4,
	r_sync_rst,
	b_full,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	b_non_empty,
	r_val,
	fifo_wr,
	src_payload,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_7;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_6;
output 	q_b_5;
output 	q_b_4;
input 	r_sync_rst;
output 	b_full;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	b_non_empty;
input 	r_val;
input 	fifo_wr;
input 	src_payload;
input 	src_payload1;
input 	src_payload2;
input 	src_payload3;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



processor_scfifo_2 wfifo(
	.q({q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.r_sync_rst(r_sync_rst),
	.b_full(b_full),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.b_non_empty(b_non_empty),
	.r_val(r_val),
	.wrreq(fifo_wr),
	.data({src_payload,src_payload5,src_payload6,src_payload7,src_payload4,src_payload3,src_payload2,src_payload1}),
	.clock(clk_clk));

endmodule

module processor_scfifo_2 (
	q,
	r_sync_rst,
	b_full,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	b_non_empty,
	r_val,
	wrreq,
	data,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	r_sync_rst;
output 	b_full;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	b_non_empty;
input 	r_val;
input 	wrreq;
input 	[7:0] data;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



processor_scfifo_cr21_1 auto_generated(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.r_sync_rst(r_sync_rst),
	.b_full(b_full),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.b_non_empty(b_non_empty),
	.r_val(r_val),
	.wrreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.clock(clock));

endmodule

module processor_scfifo_cr21_1 (
	q,
	r_sync_rst,
	b_full,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	b_non_empty,
	r_val,
	wrreq,
	data,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	r_sync_rst;
output 	b_full;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	b_non_empty;
input 	r_val;
input 	wrreq;
input 	[7:0] data;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



processor_a_dpfifo_e011_1 dpfifo(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.r_sync_rst(r_sync_rst),
	.b_full(b_full),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.b_non_empty(b_non_empty),
	.r_val(r_val),
	.wreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.clock(clock));

endmodule

module processor_a_dpfifo_e011_1 (
	q,
	r_sync_rst,
	b_full,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	b_non_empty,
	r_val,
	wreq,
	data,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	r_sync_rst;
output 	b_full;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	b_non_empty;
input 	r_val;
input 	wreq;
input 	[7:0] data;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \wr_ptr|counter_reg_bit[5]~q ;
wire \rd_ptr_count|counter_reg_bit[0]~q ;
wire \rd_ptr_count|counter_reg_bit[1]~q ;
wire \rd_ptr_count|counter_reg_bit[2]~q ;
wire \rd_ptr_count|counter_reg_bit[3]~q ;
wire \rd_ptr_count|counter_reg_bit[4]~q ;
wire \rd_ptr_count|counter_reg_bit[5]~q ;


processor_cntr_qnb_3 wr_ptr(
	.r_sync_rst(r_sync_rst),
	.fifo_wr(wreq),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\wr_ptr|counter_reg_bit[5]~q ),
	.clock(clock));

processor_cntr_qnb_2 rd_ptr_count(
	.r_sync_rst(r_sync_rst),
	.r_val(r_val),
	.counter_reg_bit_0(\rd_ptr_count|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_count|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_count|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_count|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\rd_ptr_count|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\rd_ptr_count|counter_reg_bit[5]~q ),
	.clock(clock));

processor_altsyncram_gio1_1 FIFOram(
	.q_b({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.clocken1(r_val),
	.wren_a(wreq),
	.data_a({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_a({\wr_ptr|counter_reg_bit[5]~q ,\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.address_b({\rd_ptr_count|counter_reg_bit[5]~q ,\rd_ptr_count|counter_reg_bit[4]~q ,\rd_ptr_count|counter_reg_bit[3]~q ,\rd_ptr_count|counter_reg_bit[2]~q ,\rd_ptr_count|counter_reg_bit[1]~q ,\rd_ptr_count|counter_reg_bit[0]~q }),
	.clock1(clock),
	.clock0(clock));

processor_a_fefifo_7cf_1 fifo_state(
	.r_sync_rst(r_sync_rst),
	.b_full1(b_full),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.b_non_empty1(b_non_empty),
	.r_val(r_val),
	.wreq(wreq),
	.clock(clock));

endmodule

module processor_a_fefifo_7cf_1 (
	r_sync_rst,
	b_full1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	b_non_empty1,
	r_val,
	wreq,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	b_full1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	b_non_empty1;
input 	r_val;
input 	wreq;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \_~0_combout ;
wire \b_full~0_combout ;
wire \b_full~1_combout ;
wire \b_full~2_combout ;
wire \b_non_empty~0_combout ;
wire \b_non_empty~1_combout ;
wire \b_non_empty~2_combout ;


processor_cntr_6o7_1 count_usedw(
	.r_sync_rst(r_sync_rst),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.updown(wreq),
	._(\_~0_combout ),
	.clock(clock));

cyclone10lp_lcell_comb \_~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(wreq),
	.datad(r_val),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h0FF0;
defparam \_~0 .sum_lutc_input = "datac";

dffeas b_full(
	.clk(clock),
	.d(\b_full~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_full1),
	.prn(vcc));
defparam b_full.is_wysiwyg = "true";
defparam b_full.power_up = "low";

dffeas b_non_empty(
	.clk(clock),
	.d(\b_non_empty~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_non_empty1),
	.prn(vcc));
defparam b_non_empty.is_wysiwyg = "true";
defparam b_non_empty.power_up = "low";

cyclone10lp_lcell_comb \b_full~0 (
	.dataa(counter_reg_bit_5),
	.datab(counter_reg_bit_4),
	.datac(wreq),
	.datad(b_non_empty1),
	.cin(gnd),
	.combout(\b_full~0_combout ),
	.cout());
defparam \b_full~0 .lut_mask = 16'hFFFE;
defparam \b_full~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \b_full~1 (
	.dataa(counter_reg_bit_3),
	.datab(counter_reg_bit_2),
	.datac(counter_reg_bit_1),
	.datad(counter_reg_bit_0),
	.cin(gnd),
	.combout(\b_full~1_combout ),
	.cout());
defparam \b_full~1 .lut_mask = 16'hFFFE;
defparam \b_full~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \b_full~2 (
	.dataa(b_full1),
	.datab(\b_full~0_combout ),
	.datac(\b_full~1_combout ),
	.datad(r_val),
	.cin(gnd),
	.combout(\b_full~2_combout ),
	.cout());
defparam \b_full~2 .lut_mask = 16'hFEFF;
defparam \b_full~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \b_non_empty~0 (
	.dataa(counter_reg_bit_5),
	.datab(counter_reg_bit_4),
	.datac(counter_reg_bit_2),
	.datad(counter_reg_bit_1),
	.cin(gnd),
	.combout(\b_non_empty~0_combout ),
	.cout());
defparam \b_non_empty~0 .lut_mask = 16'hFFFE;
defparam \b_non_empty~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \b_non_empty~1 (
	.dataa(counter_reg_bit_3),
	.datab(\b_non_empty~0_combout ),
	.datac(counter_reg_bit_0),
	.datad(r_val),
	.cin(gnd),
	.combout(\b_non_empty~1_combout ),
	.cout());
defparam \b_non_empty~1 .lut_mask = 16'hEFFF;
defparam \b_non_empty~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \b_non_empty~2 (
	.dataa(b_full1),
	.datab(wreq),
	.datac(b_non_empty1),
	.datad(\b_non_empty~1_combout ),
	.cin(gnd),
	.combout(\b_non_empty~2_combout ),
	.cout());
defparam \b_non_empty~2 .lut_mask = 16'hFFFE;
defparam \b_non_empty~2 .sum_lutc_input = "datac";

endmodule

module processor_cntr_6o7_1 (
	r_sync_rst,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	updown,
	_,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	updown;
input 	_;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita0~combout ;


dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

cyclone10lp_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cyclone10lp_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cyclone10lp_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cyclone10lp_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cyclone10lp_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5A6F;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cyclone10lp_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module processor_altsyncram_gio1_1 (
	q_b,
	clocken1,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_b;
input 	clocken1;
input 	wren_a;
input 	[7:0] data_a;
input 	[5:0] address_a;
input 	[5:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

cyclone10lp_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk1_core_clock_enable = "ena1";
defparam ram_block1a7.clk1_input_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "processor_jtag_uart_0:jtag_uart_0|processor_jtag_uart_0_scfifo_w:the_processor_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_cr21:auto_generated|a_dpfifo_e011:dpfifo|altsyncram_gio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 6;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 63;
defparam ram_block1a7.port_a_logical_ram_depth = 64;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 6;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 63;
defparam ram_block1a7.port_b_logical_ram_depth = 64;
defparam ram_block1a7.port_b_logical_ram_width = 8;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk1_core_clock_enable = "ena1";
defparam ram_block1a0.clk1_input_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "processor_jtag_uart_0:jtag_uart_0|processor_jtag_uart_0_scfifo_w:the_processor_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_cr21:auto_generated|a_dpfifo_e011:dpfifo|altsyncram_gio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 6;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 63;
defparam ram_block1a0.port_a_logical_ram_depth = 64;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 6;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 63;
defparam ram_block1a0.port_b_logical_ram_depth = 64;
defparam ram_block1a0.port_b_logical_ram_width = 8;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk1_core_clock_enable = "ena1";
defparam ram_block1a1.clk1_input_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "processor_jtag_uart_0:jtag_uart_0|processor_jtag_uart_0_scfifo_w:the_processor_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_cr21:auto_generated|a_dpfifo_e011:dpfifo|altsyncram_gio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 6;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 63;
defparam ram_block1a1.port_a_logical_ram_depth = 64;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 6;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 63;
defparam ram_block1a1.port_b_logical_ram_depth = 64;
defparam ram_block1a1.port_b_logical_ram_width = 8;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk1_core_clock_enable = "ena1";
defparam ram_block1a2.clk1_input_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "processor_jtag_uart_0:jtag_uart_0|processor_jtag_uart_0_scfifo_w:the_processor_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_cr21:auto_generated|a_dpfifo_e011:dpfifo|altsyncram_gio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 6;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 63;
defparam ram_block1a2.port_a_logical_ram_depth = 64;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 6;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 63;
defparam ram_block1a2.port_b_logical_ram_depth = 64;
defparam ram_block1a2.port_b_logical_ram_width = 8;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk1_core_clock_enable = "ena1";
defparam ram_block1a3.clk1_input_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "processor_jtag_uart_0:jtag_uart_0|processor_jtag_uart_0_scfifo_w:the_processor_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_cr21:auto_generated|a_dpfifo_e011:dpfifo|altsyncram_gio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 6;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 63;
defparam ram_block1a3.port_a_logical_ram_depth = 64;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 6;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 63;
defparam ram_block1a3.port_b_logical_ram_depth = 64;
defparam ram_block1a3.port_b_logical_ram_width = 8;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk1_core_clock_enable = "ena1";
defparam ram_block1a6.clk1_input_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "processor_jtag_uart_0:jtag_uart_0|processor_jtag_uart_0_scfifo_w:the_processor_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_cr21:auto_generated|a_dpfifo_e011:dpfifo|altsyncram_gio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 6;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 63;
defparam ram_block1a6.port_a_logical_ram_depth = 64;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 6;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 63;
defparam ram_block1a6.port_b_logical_ram_depth = 64;
defparam ram_block1a6.port_b_logical_ram_width = 8;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk1_core_clock_enable = "ena1";
defparam ram_block1a5.clk1_input_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "processor_jtag_uart_0:jtag_uart_0|processor_jtag_uart_0_scfifo_w:the_processor_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_cr21:auto_generated|a_dpfifo_e011:dpfifo|altsyncram_gio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 6;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 63;
defparam ram_block1a5.port_a_logical_ram_depth = 64;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 6;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 63;
defparam ram_block1a5.port_b_logical_ram_depth = 64;
defparam ram_block1a5.port_b_logical_ram_width = 8;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk1_core_clock_enable = "ena1";
defparam ram_block1a4.clk1_input_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "processor_jtag_uart_0:jtag_uart_0|processor_jtag_uart_0_scfifo_w:the_processor_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_cr21:auto_generated|a_dpfifo_e011:dpfifo|altsyncram_gio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 6;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 63;
defparam ram_block1a4.port_a_logical_ram_depth = 64;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 6;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 63;
defparam ram_block1a4.port_b_logical_ram_depth = 64;
defparam ram_block1a4.port_b_logical_ram_width = 8;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

endmodule

module processor_cntr_qnb_2 (
	r_sync_rst,
	r_val,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	r_val;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cyclone10lp_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cyclone10lp_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cyclone10lp_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cyclone10lp_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cyclone10lp_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cyclone10lp_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module processor_cntr_qnb_3 (
	r_sync_rst,
	fifo_wr,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	fifo_wr;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cyclone10lp_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cyclone10lp_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cyclone10lp_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cyclone10lp_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cyclone10lp_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cyclone10lp_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module processor_processor_LED (
	data_out_0,
	data_out_1,
	d_writedata_0,
	r_sync_rst,
	saved_grant_0,
	src_payload,
	saved_grant_1,
	src_valid,
	src_valid1,
	mem_used_1,
	always0,
	read_mux_out,
	read_mux_out1,
	wait_latency_counter_1,
	wait_latency_counter_0,
	d_writedata_1,
	readdata_0,
	readdata_1,
	clk)/* synthesis synthesis_greybox=1 */;
output 	data_out_0;
output 	data_out_1;
input 	d_writedata_0;
input 	r_sync_rst;
input 	saved_grant_0;
input 	src_payload;
input 	saved_grant_1;
input 	src_valid;
input 	src_valid1;
input 	mem_used_1;
output 	always0;
input 	read_mux_out;
input 	read_mux_out1;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	d_writedata_1;
output 	readdata_0;
output 	readdata_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \data_out[0]~0_combout ;
wire \Equal0~0_combout ;
wire \always0~1_combout ;
wire \data_out[1]~1_combout ;


dffeas \data_out[0] (
	.clk(clk),
	.d(\data_out[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_0),
	.prn(vcc));
defparam \data_out[0] .is_wysiwyg = "true";
defparam \data_out[0] .power_up = "low";

dffeas \data_out[1] (
	.clk(clk),
	.d(\data_out[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_1),
	.prn(vcc));
defparam \data_out[1] .is_wysiwyg = "true";
defparam \data_out[1] .power_up = "low";

cyclone10lp_lcell_comb \always0~0 (
	.dataa(src_payload),
	.datab(src_valid),
	.datac(src_valid1),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(always0),
	.cout());
defparam \always0~0 .lut_mask = 16'hFEFF;
defparam \always0~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(data_out_0),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(readdata_0),
	.cout());
defparam \readdata[0] .lut_mask = 16'h0FFF;
defparam \readdata[0] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(data_out_1),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(readdata_1),
	.cout());
defparam \readdata[1] .lut_mask = 16'h0FFF;
defparam \readdata[1] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \data_out[0]~0 (
	.dataa(d_writedata_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_out[0]~0_combout ),
	.cout());
defparam \data_out[0]~0 .lut_mask = 16'h5555;
defparam \data_out[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal0~0 (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(read_mux_out),
	.datad(read_mux_out1),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hEFFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \always0~1 (
	.dataa(always0),
	.datab(\Equal0~0_combout ),
	.datac(wait_latency_counter_1),
	.datad(wait_latency_counter_0),
	.cin(gnd),
	.combout(\always0~1_combout ),
	.cout());
defparam \always0~1 .lut_mask = 16'hBFFF;
defparam \always0~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \data_out[1]~1 (
	.dataa(d_writedata_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_out[1]~1_combout ),
	.cout());
defparam \data_out[1]~1 .lut_mask = 16'h5555;
defparam \data_out[1]~1 .sum_lutc_input = "datac";

endmodule

module processor_processor_mm_interconnect_0 (
	W_alu_result_7,
	W_alu_result_16,
	W_alu_result_15,
	W_alu_result_14,
	W_alu_result_13,
	W_alu_result_12,
	W_alu_result_11,
	W_alu_result_10,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_4,
	W_alu_result_5,
	W_alu_result_6,
	W_alu_result_2,
	W_alu_result_3,
	q_a_0,
	q_a_22,
	av_readdata_pre_22,
	q_a_23,
	q_a_14,
	q_a_15,
	q_a_11,
	q_a_13,
	q_a_16,
	av_readdata_pre_16,
	q_a_12,
	q_a_10,
	q_a_9,
	q_a_8,
	q_a_21,
	av_readdata_pre_21,
	q_a_20,
	av_readdata_pre_20,
	q_a_19,
	av_readdata_pre_19,
	q_a_18,
	av_readdata_pre_18,
	q_a_17,
	av_readdata_pre_17,
	readdata_0,
	d_writedata_24,
	d_writedata_25,
	d_writedata_26,
	readdata_1,
	readdata_3,
	readdata_2,
	d_writedata_27,
	d_writedata_28,
	d_writedata_29,
	d_writedata_30,
	d_writedata_31,
	d_writedata_0,
	r_sync_rst,
	saved_grant_0,
	d_write,
	src_payload,
	saved_grant_1,
	rst1,
	i_read,
	F_pc_5,
	F_pc_14,
	F_pc_13,
	F_pc_12,
	F_pc_11,
	F_pc_10,
	F_pc_9,
	F_pc_8,
	F_pc_7,
	F_pc_6,
	F_pc_2,
	F_pc_3,
	F_pc_4,
	src_valid,
	d_read,
	src_valid1,
	mem_used_1,
	always0,
	F_pc_1,
	F_pc_0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	d_writedata_1,
	saved_grant_01,
	src_payload1,
	saved_grant_11,
	src_valid2,
	src_valid3,
	mem_used_11,
	always01,
	wait_latency_counter_11,
	wait_latency_counter_01,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	saved_grant_02,
	src_payload2,
	saved_grant_12,
	src_valid4,
	src_valid5,
	mem_used_12,
	always02,
	wait_latency_counter_12,
	wait_latency_counter_02,
	src0_valid,
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	src0_valid1,
	read_latency_shift_reg_01,
	mem_74_01,
	mem_56_01,
	src0_valid2,
	src0_valid3,
	WideOr1,
	src0_valid4,
	read_latency_shift_reg_02,
	mem_74_02,
	mem_56_02,
	src0_valid5,
	src0_valid6,
	WideOr11,
	WideOr12,
	saved_grant_03,
	mem_used_13,
	mem_used_14,
	wait_latency_counter_13,
	av_waitrequest,
	mem_used_15,
	saved_grant_04,
	saved_grant_05,
	waitrequest,
	mem_used_16,
	saved_grant_06,
	saved_grant_13,
	nios2_gen2_0_data_master_waitrequest,
	src1_valid,
	src1_valid1,
	src1_valid2,
	src1_valid3,
	WideOr13,
	src1_valid4,
	src_payload3,
	src_payload4,
	WideOr14,
	uav_write,
	d_writedata_9,
	src_payload5,
	src_data_38,
	src_data_39,
	src_data_40,
	WideOr15,
	uart_0_s1_begintransfer,
	src_data_56,
	WideOr16,
	WideOr17,
	WideOr18,
	src_data_561,
	rx_rd_strobe_onset,
	rf_source_valid,
	hbreak_enabled,
	src_data_0,
	av_readdata_pre_221,
	av_readdata_pre_23,
	av_readdata_pre_24,
	av_readdata_pre_25,
	av_readdata_pre_26,
	src_data_01,
	src_data_02,
	src_data_03,
	av_readdata_pre_1,
	av_readdata_pre_11,
	av_readdata_pre_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	av_readdata_pre_15,
	av_readdata_pre_4,
	av_readdata_pre_41,
	av_readdata_pre_42,
	av_readdata_pre_43,
	av_readdata_pre_3,
	src_payload6,
	av_readdata_pre_31,
	av_readdata_pre_32,
	av_readdata_pre_33,
	av_readdata_pre_2,
	av_readdata_pre_27,
	av_readdata_pre_28,
	av_readdata_pre_29,
	av_readdata_pre_210,
	src_data_46,
	av_readdata_pre_5,
	av_readdata_pre_51,
	av_readdata_pre_52,
	av_readdata_pre_53,
	av_readdata_pre_141,
	av_readdata_pre_142,
	av_readdata_pre_151,
	av_readdata_pre_152,
	src_payload7,
	av_readdata_pre_111,
	av_readdata_pre_131,
	av_readdata_pre_132,
	av_readdata_pre_161,
	av_readdata_pre_121,
	av_readdata_pre_122,
	av_readdata_pre_10,
	av_readdata_pre_101,
	av_readdata_pre_9,
	av_readdata_pre_91,
	av_readdata_pre_92,
	av_readdata_pre_8,
	av_readdata_pre_81,
	av_readdata_pre_82,
	av_readdata_pre_7,
	av_readdata_pre_71,
	av_readdata_pre_72,
	av_readdata_pre_73,
	av_readdata_pre_6,
	av_readdata_pre_61,
	av_readdata_pre_62,
	av_readdata_pre_63,
	av_readdata_pre_211,
	av_readdata_pre_201,
	av_readdata_pre_191,
	av_readdata_pre_181,
	av_readdata_pre_171,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	b_full,
	src_data_8,
	readdata_01,
	readdata_02,
	src_payload16,
	src_data_381,
	src_data_391,
	src_data_401,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_461,
	src_data_47,
	src_data_48,
	src_data_49,
	src_data_50,
	d_byteenable_0,
	src_data_32,
	read_0,
	av_readdata_0,
	readdata_03,
	readdata_04,
	readdata_05,
	av_readdata_9,
	av_readdata_8,
	d_writedata_22,
	src_payload17,
	d_byteenable_2,
	src_data_34,
	readdata_22,
	b_full1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	readdata_23,
	d_writedata_23,
	src_payload18,
	readdata_24,
	src_payload19,
	d_byteenable_3,
	src_data_35,
	readdata_25,
	src_payload20,
	readdata_26,
	src_payload21,
	av_readdata_1,
	src_payload22,
	readdata_11,
	readdata_12,
	readdata_13,
	readdata_14,
	src_payload23,
	readdata_4,
	readdata_41,
	readdata_42,
	av_readdata_4,
	av_readdata_3,
	src_payload24,
	readdata_31,
	readdata_32,
	av_readdata_2,
	readdata_21,
	src_payload25,
	readdata_27,
	readdata_28,
	src_payload26,
	readdata_5,
	readdata_51,
	readdata_52,
	av_readdata_5,
	d_writedata_14,
	src_payload27,
	d_byteenable_1,
	src_data_33,
	readdata_141,
	woverflow,
	d_writedata_15,
	src_payload28,
	readdata_15,
	rvalid,
	d_writedata_11,
	src_payload29,
	readdata_111,
	d_writedata_13,
	src_payload30,
	readdata_131,
	d_writedata_16,
	src_payload31,
	readdata_16,
	counter_reg_bit_01,
	d_writedata_12,
	src_payload32,
	readdata_121,
	b_non_empty,
	av_readdata_pre_271,
	av_readdata_pre_281,
	av_readdata_pre_291,
	av_readdata_pre_30,
	av_readdata_pre_311,
	d_writedata_10,
	src_payload33,
	readdata_10,
	ac,
	readdata_9,
	readdata_91,
	src_payload34,
	readdata_8,
	readdata_81,
	d_writedata_8,
	src_payload35,
	readdata_7,
	av_readdata_7,
	src_payload36,
	readdata_71,
	readdata_72,
	readdata_6,
	av_readdata_6,
	src_payload37,
	readdata_61,
	readdata_62,
	src_payload38,
	d_writedata_21,
	src_payload39,
	readdata_211,
	counter_reg_bit_51,
	d_writedata_20,
	src_payload40,
	readdata_20,
	counter_reg_bit_41,
	src_payload41,
	d_writedata_19,
	src_payload42,
	readdata_19,
	counter_reg_bit_31,
	src_payload43,
	d_writedata_18,
	src_payload44,
	counter_reg_bit_21,
	readdata_18,
	src_payload45,
	d_writedata_17,
	src_payload46,
	counter_reg_bit_11,
	readdata_17,
	src_payload47,
	src_payload48,
	src_payload49,
	src_data_9,
	end_begintransfer,
	src_data_382,
	src_payload50,
	src_payload51,
	src_payload52,
	src_data_383,
	src_data_392,
	src_data_402,
	src_data_411,
	src_data_421,
	src_data_431,
	src_data_441,
	src_data_451,
	src_data_321,
	src_payload53,
	src_payload54,
	readdata_271,
	src_payload55,
	readdata_281,
	src_payload56,
	readdata_29,
	src_payload57,
	readdata_30,
	src_payload58,
	readdata_311,
	src_payload59,
	src_payload60,
	src_payload61,
	src_payload62,
	src_payload63,
	src_payload64,
	src_payload65,
	src_payload66,
	src_payload67,
	src_payload68,
	src_payload69,
	src_payload70,
	src_payload71,
	src_data_341,
	src_payload72,
	src_payload73,
	src_data_351,
	src_payload74,
	src_payload75,
	src_payload76,
	src_payload77,
	src_payload78,
	src_data_331,
	src_payload79,
	src_payload80,
	src_payload81,
	src_payload82,
	src_payload83,
	src_payload84,
	src_payload85,
	src_payload86,
	src_payload87,
	src_payload88,
	src_payload89,
	src_payload90,
	src_payload91,
	src_payload92,
	src_payload93,
	src_payload94,
	src_payload95,
	src_payload96,
	src_payload97,
	src_payload98,
	src_payload99,
	src_payload100,
	src_payload101,
	src_payload102,
	src_payload103,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_7;
input 	W_alu_result_16;
input 	W_alu_result_15;
input 	W_alu_result_14;
input 	W_alu_result_13;
input 	W_alu_result_12;
input 	W_alu_result_11;
input 	W_alu_result_10;
input 	W_alu_result_9;
input 	W_alu_result_8;
input 	W_alu_result_4;
input 	W_alu_result_5;
input 	W_alu_result_6;
input 	W_alu_result_2;
input 	W_alu_result_3;
input 	q_a_0;
input 	q_a_22;
output 	av_readdata_pre_22;
input 	q_a_23;
input 	q_a_14;
input 	q_a_15;
input 	q_a_11;
input 	q_a_13;
input 	q_a_16;
output 	av_readdata_pre_16;
input 	q_a_12;
input 	q_a_10;
input 	q_a_9;
input 	q_a_8;
input 	q_a_21;
output 	av_readdata_pre_21;
input 	q_a_20;
output 	av_readdata_pre_20;
input 	q_a_19;
output 	av_readdata_pre_19;
input 	q_a_18;
output 	av_readdata_pre_18;
input 	q_a_17;
output 	av_readdata_pre_17;
input 	readdata_0;
input 	d_writedata_24;
input 	d_writedata_25;
input 	d_writedata_26;
input 	readdata_1;
input 	readdata_3;
input 	readdata_2;
input 	d_writedata_27;
input 	d_writedata_28;
input 	d_writedata_29;
input 	d_writedata_30;
input 	d_writedata_31;
input 	d_writedata_0;
input 	r_sync_rst;
output 	saved_grant_0;
input 	d_write;
output 	src_payload;
output 	saved_grant_1;
input 	rst1;
input 	i_read;
input 	F_pc_5;
input 	F_pc_14;
input 	F_pc_13;
input 	F_pc_12;
input 	F_pc_11;
input 	F_pc_10;
input 	F_pc_9;
input 	F_pc_8;
input 	F_pc_7;
input 	F_pc_6;
input 	F_pc_2;
input 	F_pc_3;
input 	F_pc_4;
output 	src_valid;
input 	d_read;
output 	src_valid1;
output 	mem_used_1;
input 	always0;
input 	F_pc_1;
input 	F_pc_0;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
input 	d_writedata_1;
output 	saved_grant_01;
output 	src_payload1;
output 	saved_grant_11;
output 	src_valid2;
output 	src_valid3;
output 	mem_used_11;
input 	always01;
output 	wait_latency_counter_11;
output 	wait_latency_counter_01;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
output 	saved_grant_02;
output 	src_payload2;
output 	saved_grant_12;
output 	src_valid4;
output 	src_valid5;
output 	mem_used_12;
input 	always02;
output 	wait_latency_counter_12;
output 	wait_latency_counter_02;
output 	src0_valid;
output 	read_latency_shift_reg_0;
output 	mem_74_0;
output 	mem_56_0;
output 	src0_valid1;
output 	read_latency_shift_reg_01;
output 	mem_74_01;
output 	mem_56_01;
output 	src0_valid2;
output 	src0_valid3;
output 	WideOr1;
output 	src0_valid4;
output 	read_latency_shift_reg_02;
output 	mem_74_02;
output 	mem_56_02;
output 	src0_valid5;
output 	src0_valid6;
output 	WideOr11;
output 	WideOr12;
output 	saved_grant_03;
output 	mem_used_13;
output 	mem_used_14;
output 	wait_latency_counter_13;
input 	av_waitrequest;
output 	mem_used_15;
output 	saved_grant_04;
output 	saved_grant_05;
input 	waitrequest;
output 	mem_used_16;
output 	saved_grant_06;
output 	saved_grant_13;
output 	nios2_gen2_0_data_master_waitrequest;
output 	src1_valid;
output 	src1_valid1;
output 	src1_valid2;
output 	src1_valid3;
output 	WideOr13;
output 	src1_valid4;
output 	src_payload3;
output 	src_payload4;
output 	WideOr14;
output 	uav_write;
input 	d_writedata_9;
output 	src_payload5;
output 	src_data_38;
output 	src_data_39;
output 	src_data_40;
output 	WideOr15;
output 	uart_0_s1_begintransfer;
output 	src_data_56;
output 	WideOr16;
output 	WideOr17;
output 	WideOr18;
output 	src_data_561;
input 	rx_rd_strobe_onset;
output 	rf_source_valid;
input 	hbreak_enabled;
output 	src_data_0;
output 	av_readdata_pre_221;
output 	av_readdata_pre_23;
output 	av_readdata_pre_24;
output 	av_readdata_pre_25;
output 	av_readdata_pre_26;
output 	src_data_01;
output 	src_data_02;
output 	src_data_03;
output 	av_readdata_pre_1;
output 	av_readdata_pre_11;
output 	av_readdata_pre_12;
output 	av_readdata_pre_13;
output 	av_readdata_pre_14;
output 	av_readdata_pre_15;
output 	av_readdata_pre_4;
output 	av_readdata_pre_41;
output 	av_readdata_pre_42;
output 	av_readdata_pre_43;
output 	av_readdata_pre_3;
output 	src_payload6;
output 	av_readdata_pre_31;
output 	av_readdata_pre_32;
output 	av_readdata_pre_33;
output 	av_readdata_pre_2;
output 	av_readdata_pre_27;
output 	av_readdata_pre_28;
output 	av_readdata_pre_29;
output 	av_readdata_pre_210;
output 	src_data_46;
output 	av_readdata_pre_5;
output 	av_readdata_pre_51;
output 	av_readdata_pre_52;
output 	av_readdata_pre_53;
output 	av_readdata_pre_141;
output 	av_readdata_pre_142;
output 	av_readdata_pre_151;
output 	av_readdata_pre_152;
output 	src_payload7;
output 	av_readdata_pre_111;
output 	av_readdata_pre_131;
output 	av_readdata_pre_132;
output 	av_readdata_pre_161;
output 	av_readdata_pre_121;
output 	av_readdata_pre_122;
output 	av_readdata_pre_10;
output 	av_readdata_pre_101;
output 	av_readdata_pre_9;
output 	av_readdata_pre_91;
output 	av_readdata_pre_92;
output 	av_readdata_pre_8;
output 	av_readdata_pre_81;
output 	av_readdata_pre_82;
output 	av_readdata_pre_7;
output 	av_readdata_pre_71;
output 	av_readdata_pre_72;
output 	av_readdata_pre_73;
output 	av_readdata_pre_6;
output 	av_readdata_pre_61;
output 	av_readdata_pre_62;
output 	av_readdata_pre_63;
output 	av_readdata_pre_211;
output 	av_readdata_pre_201;
output 	av_readdata_pre_191;
output 	av_readdata_pre_181;
output 	av_readdata_pre_171;
output 	src_payload8;
output 	src_payload9;
output 	src_payload10;
output 	src_payload11;
output 	src_payload12;
output 	src_payload13;
output 	src_payload14;
output 	src_payload15;
input 	b_full;
output 	src_data_8;
input 	readdata_01;
input 	readdata_02;
output 	src_payload16;
output 	src_data_381;
output 	src_data_391;
output 	src_data_401;
output 	src_data_41;
output 	src_data_42;
output 	src_data_43;
output 	src_data_44;
output 	src_data_45;
output 	src_data_461;
output 	src_data_47;
output 	src_data_48;
output 	src_data_49;
output 	src_data_50;
input 	d_byteenable_0;
output 	src_data_32;
input 	read_0;
input 	av_readdata_0;
input 	readdata_03;
input 	readdata_04;
input 	readdata_05;
input 	av_readdata_9;
input 	av_readdata_8;
input 	d_writedata_22;
output 	src_payload17;
input 	d_byteenable_2;
output 	src_data_34;
input 	readdata_22;
input 	b_full1;
input 	counter_reg_bit_5;
input 	counter_reg_bit_4;
input 	counter_reg_bit_3;
input 	counter_reg_bit_2;
input 	counter_reg_bit_1;
input 	counter_reg_bit_0;
input 	readdata_23;
input 	d_writedata_23;
output 	src_payload18;
input 	readdata_24;
output 	src_payload19;
input 	d_byteenable_3;
output 	src_data_35;
input 	readdata_25;
output 	src_payload20;
input 	readdata_26;
output 	src_payload21;
input 	av_readdata_1;
output 	src_payload22;
input 	readdata_11;
input 	readdata_12;
input 	readdata_13;
input 	readdata_14;
output 	src_payload23;
input 	readdata_4;
input 	readdata_41;
input 	readdata_42;
input 	av_readdata_4;
input 	av_readdata_3;
output 	src_payload24;
input 	readdata_31;
input 	readdata_32;
input 	av_readdata_2;
input 	readdata_21;
output 	src_payload25;
input 	readdata_27;
input 	readdata_28;
output 	src_payload26;
input 	readdata_5;
input 	readdata_51;
input 	readdata_52;
input 	av_readdata_5;
input 	d_writedata_14;
output 	src_payload27;
input 	d_byteenable_1;
output 	src_data_33;
input 	readdata_141;
input 	woverflow;
input 	d_writedata_15;
output 	src_payload28;
input 	readdata_15;
input 	rvalid;
input 	d_writedata_11;
output 	src_payload29;
input 	readdata_111;
input 	d_writedata_13;
output 	src_payload30;
input 	readdata_131;
input 	d_writedata_16;
output 	src_payload31;
input 	readdata_16;
input 	counter_reg_bit_01;
input 	d_writedata_12;
output 	src_payload32;
input 	readdata_121;
input 	b_non_empty;
output 	av_readdata_pre_271;
output 	av_readdata_pre_281;
output 	av_readdata_pre_291;
output 	av_readdata_pre_30;
output 	av_readdata_pre_311;
input 	d_writedata_10;
output 	src_payload33;
input 	readdata_10;
input 	ac;
input 	readdata_9;
input 	readdata_91;
output 	src_payload34;
input 	readdata_8;
input 	readdata_81;
input 	d_writedata_8;
output 	src_payload35;
input 	readdata_7;
input 	av_readdata_7;
output 	src_payload36;
input 	readdata_71;
input 	readdata_72;
input 	readdata_6;
input 	av_readdata_6;
output 	src_payload37;
input 	readdata_61;
input 	readdata_62;
output 	src_payload38;
input 	d_writedata_21;
output 	src_payload39;
input 	readdata_211;
input 	counter_reg_bit_51;
input 	d_writedata_20;
output 	src_payload40;
input 	readdata_20;
input 	counter_reg_bit_41;
output 	src_payload41;
input 	d_writedata_19;
output 	src_payload42;
input 	readdata_19;
input 	counter_reg_bit_31;
output 	src_payload43;
input 	d_writedata_18;
output 	src_payload44;
input 	counter_reg_bit_21;
input 	readdata_18;
output 	src_payload45;
input 	d_writedata_17;
output 	src_payload46;
input 	counter_reg_bit_11;
input 	readdata_17;
output 	src_payload47;
output 	src_payload48;
output 	src_payload49;
output 	src_data_9;
output 	end_begintransfer;
output 	src_data_382;
output 	src_payload50;
output 	src_payload51;
output 	src_payload52;
output 	src_data_383;
output 	src_data_392;
output 	src_data_402;
output 	src_data_411;
output 	src_data_421;
output 	src_data_431;
output 	src_data_441;
output 	src_data_451;
output 	src_data_321;
output 	src_payload53;
output 	src_payload54;
input 	readdata_271;
output 	src_payload55;
input 	readdata_281;
output 	src_payload56;
input 	readdata_29;
output 	src_payload57;
input 	readdata_30;
output 	src_payload58;
input 	readdata_311;
output 	src_payload59;
output 	src_payload60;
output 	src_payload61;
output 	src_payload62;
output 	src_payload63;
output 	src_payload64;
output 	src_payload65;
output 	src_payload66;
output 	src_payload67;
output 	src_payload68;
output 	src_payload69;
output 	src_payload70;
output 	src_payload71;
output 	src_data_341;
output 	src_payload72;
output 	src_payload73;
output 	src_data_351;
output 	src_payload74;
output 	src_payload75;
output 	src_payload76;
output 	src_payload77;
output 	src_payload78;
output 	src_data_331;
output 	src_payload79;
output 	src_payload80;
output 	src_payload81;
output 	src_payload82;
output 	src_payload83;
output 	src_payload84;
output 	src_payload85;
output 	src_payload86;
output 	src_payload87;
output 	src_payload88;
output 	src_payload89;
output 	src_payload90;
output 	src_payload91;
output 	src_payload92;
output 	src_payload93;
output 	src_payload94;
output 	src_payload95;
output 	src_payload96;
output 	src_payload97;
output 	src_payload98;
output 	src_payload99;
output 	src_payload100;
output 	src_payload101;
output 	src_payload102;
output 	src_payload103;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \nios2_gen2_0_data_master_translator|write_accepted~q ;
wire \nios2_gen2_0_instruction_master_translator|read_accepted~q ;
wire \nios2_gen2_0_instruction_master_agent|cp_valid~combout ;
wire \router_001|Equal1~0_combout ;
wire \router_001|Equal4~0_combout ;
wire \router|Equal4~0_combout ;
wire \nios2_gen2_0_data_master_translator|read_accepted~q ;
wire \nios2_gen2_0_data_master_agent|cp_valid~0_combout ;
wire \router_001|Equal4~2_combout ;
wire \router|Equal6~1_combout ;
wire \nios2_gen2_0_data_master_agent|cp_valid~1_combout ;
wire \nios2_gen2_0_instruction_master_translator|uav_read~combout ;
wire \router_001|Equal6~1_combout ;
wire \led_s1_agent|cp_ready~0_combout ;
wire \jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ;
wire \jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo|mem[0][74]~q ;
wire \jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo|mem[0][56]~q ;
wire \led_s1_translator|read_latency_shift_reg[0]~q ;
wire \led_s1_agent_rsp_fifo|mem[0][74]~q ;
wire \led_s1_agent_rsp_fifo|mem[0][56]~q ;
wire \seg_en_s1_translator|read_latency_shift_reg[0]~q ;
wire \seg_en_s1_agent_rsp_fifo|mem[0][74]~q ;
wire \seg_en_s1_agent_rsp_fifo|mem[0][56]~q ;
wire \sw_s1_translator|read_latency_shift_reg[0]~q ;
wire \sw_s1_agent_rsp_fifo|mem[0][74]~q ;
wire \sw_s1_agent_rsp_fifo|mem[0][56]~q ;
wire \rsp_demux_006|src0_valid~0_combout ;
wire \uart_0_s1_translator|read_latency_shift_reg[0]~q ;
wire \uart_0_s1_agent_rsp_fifo|mem[0][74]~q ;
wire \uart_0_s1_agent_rsp_fifo|mem[0][56]~q ;
wire \router|Equal5~1_combout ;
wire \seg_en_s1_agent|cp_ready~0_combout ;
wire \router|Equal1~1_combout ;
wire \router|Equal7~0_combout ;
wire \router|Equal2~2_combout ;
wire \router|always1~0_combout ;
wire \router|always1~1_combout ;
wire \cmd_mux_007|saved_grant[0]~q ;
wire \uart_0_s1_translator|uav_waitrequest~0_combout ;
wire \cmd_demux|sink_ready~4_combout ;
wire \router|Equal4~1_combout ;
wire \seg_s1_agent|cp_ready~0_combout ;
wire \sw_s1_translator|wait_latency_counter[0]~q ;
wire \router_001|always1~0_combout ;
wire \cmd_mux_006|src_valid~2_combout ;
wire \cmd_mux_006|src_valid~4_combout ;
wire \sw_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \sw_s1_agent|m0_write~1_combout ;
wire \sw_s1_translator|wait_latency_counter[1]~q ;
wire \sw_s1_agent|cp_ready~0_combout ;
wire \cmd_demux|WideOr0~2_combout ;
wire \router_001|Equal7~0_combout ;
wire \cmd_mux|saved_grant[1]~q ;
wire \cmd_mux_001|saved_grant[1]~q ;
wire \nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|write~0_combout ;
wire \router_001|Equal1~1_combout ;
wire \cmd_mux_002|saved_grant[1]~q ;
wire \router_001|src_channel[2]~0_combout ;
wire \router_001|Equal2~2_combout ;
wire \router_001|src_channel[2]~1_combout ;
wire \router_001|src_channel[2]~2_combout ;
wire \cmd_mux_007|saved_grant[1]~q ;
wire \router_001|Equal5~1_combout ;
wire \seg_en_s1_agent|cp_ready~2_combout ;
wire \router_001|Equal4~3_combout ;
wire \router_001|always1~1_combout ;
wire \sw_s1_agent|cp_ready~combout ;
wire \cmd_mux_003|WideOr1~combout ;
wire \nios2_gen2_0_data_master_translator|uav_read~combout ;
wire \cmd_mux_003|src_data[56]~combout ;
wire \cmd_demux_001|src5_valid~0_combout ;
wire \seg_s1_agent_rsp_fifo|write~1_combout ;
wire \cmd_mux_005|WideOr1~combout ;
wire \cmd_mux_005|src_data[56]~combout ;
wire \cmd_mux_004|WideOr1~combout ;
wire \cmd_mux_004|src_data[56]~combout ;
wire \cmd_demux_001|src0_valid~0_combout ;
wire \cmd_demux_001|src1_valid~0_combout ;
wire \nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|mem~0_combout ;
wire \cmd_demux|src2_valid~2_combout ;
wire \cmd_demux_001|src2_valid~0_combout ;
wire \onchip_memory2_0_s1_agent_rsp_fifo|mem~0_combout ;
wire \onchip_memory2_0_s1_translator|read_latency_shift_reg~0_combout ;
wire \led_s1_translator|read_latency_shift_reg~0_combout ;
wire \cmd_mux_006|WideOr1~combout ;
wire \cmd_mux_006|src_data[56]~combout ;
wire \uart_0_s1_translator|read_latency_shift_reg~0_combout ;
wire \cmd_demux_001|src6_valid~0_combout ;
wire \sw_s1_translator|read_latency_shift_reg~1_combout ;
wire \seg_s1_translator|av_readdata_pre[0]~q ;
wire \seg_en_s1_translator|av_readdata_pre[0]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[0]~q ;
wire \nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[0]~q ;
wire \uart_0_s1_translator|av_readdata_pre[0]~q ;
wire \led_s1_translator|av_readdata_pre[0]~q ;
wire \sw_s1_translator|av_readdata_pre[0]~q ;
wire \cmd_demux_001|src3_valid~2_combout ;
wire \cmd_mux_004|src_valid~6_combout ;
wire \cmd_demux_001|src4_valid~2_combout ;
wire \cmd_demux_001|src7_valid~2_combout ;


processor_processor_mm_interconnect_0_router_1 router_001(
	.i_read(i_read),
	.read_accepted(\nios2_gen2_0_instruction_master_translator|read_accepted~q ),
	.F_pc_5(F_pc_5),
	.F_pc_14(F_pc_14),
	.F_pc_13(F_pc_13),
	.F_pc_12(F_pc_12),
	.F_pc_11(F_pc_11),
	.Equal1(\router_001|Equal1~0_combout ),
	.F_pc_10(F_pc_10),
	.F_pc_9(F_pc_9),
	.F_pc_8(F_pc_8),
	.F_pc_7(F_pc_7),
	.F_pc_6(F_pc_6),
	.Equal4(\router_001|Equal4~0_combout ),
	.F_pc_2(F_pc_2),
	.F_pc_3(F_pc_3),
	.F_pc_4(F_pc_4),
	.F_pc_1(F_pc_1),
	.Equal41(\router_001|Equal4~2_combout ),
	.Equal6(\router_001|Equal6~1_combout ),
	.always1(\router_001|always1~0_combout ),
	.Equal7(\router_001|Equal7~0_combout ),
	.Equal11(\router_001|Equal1~1_combout ),
	.src_channel_2(\router_001|src_channel[2]~0_combout ),
	.Equal2(\router_001|Equal2~2_combout ),
	.src_channel_21(\router_001|src_channel[2]~1_combout ),
	.src_channel_22(\router_001|src_channel[2]~2_combout ),
	.Equal5(\router_001|Equal5~1_combout ),
	.Equal42(\router_001|Equal4~3_combout ),
	.always11(\router_001|always1~1_combout ));

processor_processor_mm_interconnect_0_router router(
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_16(W_alu_result_16),
	.W_alu_result_15(W_alu_result_15),
	.W_alu_result_14(W_alu_result_14),
	.W_alu_result_13(W_alu_result_13),
	.W_alu_result_12(W_alu_result_12),
	.W_alu_result_11(W_alu_result_11),
	.W_alu_result_10(W_alu_result_10),
	.W_alu_result_9(W_alu_result_9),
	.W_alu_result_8(W_alu_result_8),
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_6(W_alu_result_6),
	.W_alu_result_3(W_alu_result_3),
	.Equal4(\router|Equal4~0_combout ),
	.read_accepted(\nios2_gen2_0_data_master_translator|read_accepted~q ),
	.d_read(d_read),
	.Equal6(\router|Equal6~1_combout ),
	.Equal5(\router|Equal5~1_combout ),
	.Equal1(\router|Equal1~1_combout ),
	.Equal7(\router|Equal7~0_combout ),
	.Equal2(\router|Equal2~2_combout ),
	.always1(\router|always1~0_combout ),
	.always11(\router|always1~1_combout ),
	.Equal41(\router|Equal4~1_combout ));

processor_altera_avalon_sc_fifo_7 uart_0_s1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.read_latency_shift_reg_0(\uart_0_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\uart_0_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\uart_0_s1_agent_rsp_fifo|mem[0][56]~q ),
	.mem_used_1(mem_used_14),
	.uav_waitrequest(\uart_0_s1_translator|uav_waitrequest~0_combout ),
	.saved_grant_1(\cmd_mux_007|saved_grant[1]~q ),
	.WideOr1(WideOr15),
	.src_data_56(src_data_561),
	.read_latency_shift_reg(\uart_0_s1_translator|read_latency_shift_reg~0_combout ),
	.clk(clk_clk));

processor_altera_avalon_sc_fifo_6 sw_s1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.read_latency_shift_reg_0(\sw_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\sw_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\sw_s1_agent_rsp_fifo|mem[0][56]~q ),
	.saved_grant_1(saved_grant_13),
	.mem_used_1(\sw_s1_agent_rsp_fifo|mem_used[1]~q ),
	.cp_ready(\sw_s1_agent|cp_ready~0_combout ),
	.cp_ready1(\sw_s1_agent|cp_ready~combout ),
	.WideOr1(\cmd_mux_006|WideOr1~combout ),
	.src_data_56(\cmd_mux_006|src_data[56]~combout ),
	.read_latency_shift_reg(\sw_s1_translator|read_latency_shift_reg~1_combout ),
	.clk(clk_clk));

processor_altera_merlin_slave_agent_6 sw_s1_agent(
	.d_write(d_write),
	.write_accepted(\nios2_gen2_0_data_master_translator|write_accepted~q ),
	.rst1(rst1),
	.saved_grant_0(saved_grant_06),
	.wait_latency_counter_0(\sw_s1_translator|wait_latency_counter[0]~q ),
	.src_valid(\cmd_mux_006|src_valid~2_combout ),
	.src_valid1(\cmd_mux_006|src_valid~4_combout ),
	.mem_used_1(\sw_s1_agent_rsp_fifo|mem_used[1]~q ),
	.m0_write(\sw_s1_agent|m0_write~1_combout ),
	.wait_latency_counter_1(\sw_s1_translator|wait_latency_counter[1]~q ),
	.cp_ready1(\sw_s1_agent|cp_ready~0_combout ),
	.cp_ready2(\sw_s1_agent|cp_ready~combout ));

processor_altera_avalon_sc_fifo_5 seg_s1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.rst1(rst1),
	.saved_grant_1(saved_grant_11),
	.src_valid(src_valid2),
	.src_valid1(src_valid3),
	.mem_used_1(mem_used_11),
	.always0(always01),
	.wait_latency_counter_1(wait_latency_counter_11),
	.wait_latency_counter_0(wait_latency_counter_01),
	.read_latency_shift_reg_0(read_latency_shift_reg_02),
	.mem_74_0(mem_74_02),
	.mem_56_0(mem_56_02),
	.cp_ready(\seg_s1_agent|cp_ready~0_combout ),
	.write(\seg_s1_agent_rsp_fifo|write~1_combout ),
	.WideOr1(\cmd_mux_005|WideOr1~combout ),
	.src_data_56(\cmd_mux_005|src_data[56]~combout ),
	.clk(clk_clk));

processor_altera_merlin_slave_agent_5 seg_s1_agent(
	.rst1(rst1),
	.always0(always01),
	.wait_latency_counter_1(wait_latency_counter_11),
	.wait_latency_counter_0(wait_latency_counter_01),
	.cp_ready(\seg_s1_agent|cp_ready~0_combout ));

processor_altera_avalon_sc_fifo_4 seg_en_s1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.saved_grant_0(saved_grant_02),
	.saved_grant_1(saved_grant_12),
	.src_valid(src_valid4),
	.mem_used_1(mem_used_12),
	.read_latency_shift_reg_0(\seg_en_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\seg_en_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\seg_en_s1_agent_rsp_fifo|mem[0][56]~q ),
	.cp_ready(\seg_en_s1_agent|cp_ready~0_combout ),
	.src_data_56(\cmd_mux_004|src_data[56]~combout ),
	.src_valid1(\cmd_mux_004|src_valid~6_combout ),
	.clk(clk_clk));

processor_altera_merlin_slave_agent_4 seg_en_s1_agent(
	.rst1(rst1),
	.mem_used_1(mem_used_12),
	.always0(always02),
	.wait_latency_counter_1(wait_latency_counter_12),
	.wait_latency_counter_0(wait_latency_counter_02),
	.cp_ready(\seg_en_s1_agent|cp_ready~0_combout ),
	.cp_ready1(\seg_en_s1_agent|cp_ready~2_combout ));

processor_altera_avalon_sc_fifo_1 led_s1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.saved_grant_1(saved_grant_1),
	.mem_used_1(mem_used_1),
	.cp_ready(\led_s1_agent|cp_ready~0_combout ),
	.read_latency_shift_reg_0(\led_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\led_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\led_s1_agent_rsp_fifo|mem[0][56]~q ),
	.WideOr1(\cmd_mux_003|WideOr1~combout ),
	.src_data_56(\cmd_mux_003|src_data[56]~combout ),
	.read_latency_shift_reg(\led_s1_translator|read_latency_shift_reg~0_combout ),
	.clk(clk_clk));

processor_altera_merlin_slave_agent_1 led_s1_agent(
	.rst1(rst1),
	.always0(always0),
	.wait_latency_counter_1(wait_latency_counter_1),
	.wait_latency_counter_0(wait_latency_counter_0),
	.cp_ready(\led_s1_agent|cp_ready~0_combout ));

processor_altera_avalon_sc_fifo_3 onchip_memory2_0_s1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.rst1(rst1),
	.uav_read(\nios2_gen2_0_instruction_master_translator|uav_read~combout ),
	.read_latency_shift_reg_0(read_latency_shift_reg_01),
	.mem_74_0(mem_74_01),
	.mem_56_0(mem_56_01),
	.saved_grant_0(saved_grant_03),
	.mem_used_1(mem_used_13),
	.saved_grant_1(\cmd_mux_002|saved_grant[1]~q ),
	.uav_read1(\nios2_gen2_0_data_master_translator|uav_read~combout ),
	.WideOr1(WideOr18),
	.mem(\onchip_memory2_0_s1_agent_rsp_fifo|mem~0_combout ),
	.read_latency_shift_reg(\onchip_memory2_0_s1_translator|read_latency_shift_reg~0_combout ),
	.clk(clk_clk));

processor_altera_avalon_sc_fifo_2 nios2_gen2_0_debug_mem_slave_agent_rsp_fifo(
	.reset(r_sync_rst),
	.uav_read(\nios2_gen2_0_instruction_master_translator|uav_read~combout ),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.mem_74_0(mem_74_0),
	.mem_56_0(mem_56_0),
	.saved_grant_0(saved_grant_05),
	.waitrequest(waitrequest),
	.mem_used_1(mem_used_16),
	.saved_grant_1(\cmd_mux_001|saved_grant[1]~q ),
	.write(\nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|write~0_combout ),
	.uav_read1(\nios2_gen2_0_data_master_translator|uav_read~combout ),
	.WideOr1(WideOr17),
	.mem(\nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|mem~0_combout ),
	.rf_source_valid(rf_source_valid),
	.clk(clk_clk));

processor_altera_merlin_slave_agent_2 nios2_gen2_0_debug_mem_slave_agent(
	.WideOr1(WideOr17),
	.mem(\nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|mem~0_combout ),
	.rf_source_valid(rf_source_valid));

processor_altera_avalon_sc_fifo jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo(
	.reset(r_sync_rst),
	.read_latency_shift_reg_0(\jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo|mem[0][56]~q ),
	.av_waitrequest(av_waitrequest),
	.mem_used_1(mem_used_15),
	.sink_ready(\cmd_demux|sink_ready~4_combout ),
	.saved_grant_1(\cmd_mux|saved_grant[1]~q ),
	.src_data_56(src_data_56),
	.WideOr1(WideOr16),
	.clk(clk_clk));

processor_altera_merlin_master_agent_1 nios2_gen2_0_instruction_master_agent(
	.rst1(rst1),
	.i_read(i_read),
	.read_accepted(\nios2_gen2_0_instruction_master_translator|read_accepted~q ),
	.cp_valid1(\nios2_gen2_0_instruction_master_agent|cp_valid~combout ));

processor_altera_merlin_master_agent nios2_gen2_0_data_master_agent(
	.d_write(d_write),
	.write_accepted(\nios2_gen2_0_data_master_translator|write_accepted~q ),
	.rst1(rst1),
	.read_accepted(\nios2_gen2_0_data_master_translator|read_accepted~q ),
	.d_read(d_read),
	.cp_valid(\nios2_gen2_0_data_master_agent|cp_valid~0_combout ),
	.cp_valid1(\nios2_gen2_0_data_master_agent|cp_valid~1_combout ));

processor_altera_merlin_slave_translator_7 uart_0_s1_translator(
	.reset(r_sync_rst),
	.d_write(d_write),
	.write_accepted(\nios2_gen2_0_data_master_translator|write_accepted~q ),
	.rst1(rst1),
	.read_latency_shift_reg_0(\uart_0_s1_translator|read_latency_shift_reg[0]~q ),
	.saved_grant_0(\cmd_mux_007|saved_grant[0]~q ),
	.mem_used_1(mem_used_14),
	.wait_latency_counter_1(wait_latency_counter_13),
	.uav_waitrequest(\uart_0_s1_translator|uav_waitrequest~0_combout ),
	.WideOr1(WideOr15),
	.av_begintransfer(uart_0_s1_begintransfer),
	.src_data_56(src_data_561),
	.read_latency_shift_reg(\uart_0_s1_translator|read_latency_shift_reg~0_combout ),
	.rx_rd_strobe_onset(rx_rd_strobe_onset),
	.av_readdata_pre_0(\uart_0_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(av_readdata_pre_12),
	.av_readdata_pre_4(av_readdata_pre_41),
	.av_readdata_pre_3(av_readdata_pre_32),
	.av_readdata_pre_2(av_readdata_pre_210),
	.av_readdata_pre_5(av_readdata_pre_51),
	.av_readdata_pre_9(av_readdata_pre_92),
	.av_readdata_pre_8(av_readdata_pre_82),
	.av_readdata_pre_7(av_readdata_pre_73),
	.av_readdata_pre_6(av_readdata_pre_63),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_91,readdata_81,readdata_72,readdata_62,readdata_51,readdata_41,readdata_31,readdata_28,readdata_11,readdata_03}),
	.end_begintransfer1(end_begintransfer),
	.clk(clk_clk));

processor_altera_merlin_slave_translator_6 sw_s1_translator(
	.reset(r_sync_rst),
	.rst1(rst1),
	.read_latency_shift_reg_0(\sw_s1_translator|read_latency_shift_reg[0]~q ),
	.saved_grant_0(saved_grant_06),
	.wait_latency_counter_0(\sw_s1_translator|wait_latency_counter[0]~q ),
	.src_valid(\cmd_mux_006|src_valid~2_combout ),
	.src_valid1(\cmd_mux_006|src_valid~4_combout ),
	.mem_used_1(\sw_s1_agent_rsp_fifo|mem_used[1]~q ),
	.m0_write(\sw_s1_agent|m0_write~1_combout ),
	.wait_latency_counter_1(\sw_s1_translator|wait_latency_counter[1]~q ),
	.cp_ready(\sw_s1_agent|cp_ready~0_combout ),
	.uav_write(uav_write),
	.WideOr1(\cmd_mux_006|WideOr1~combout ),
	.src_data_56(\cmd_mux_006|src_data[56]~combout ),
	.read_latency_shift_reg(\sw_s1_translator|read_latency_shift_reg~1_combout ),
	.av_readdata_pre_0(\sw_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_05}),
	.clk(clk_clk));

processor_altera_merlin_slave_translator_5 seg_s1_translator(
	.reset(r_sync_rst),
	.rst1(rst1),
	.saved_grant_0(saved_grant_01),
	.src_valid(src_valid2),
	.src_valid1(src_valid3),
	.mem_used_1(mem_used_11),
	.always0(always01),
	.wait_latency_counter_1(wait_latency_counter_11),
	.wait_latency_counter_0(wait_latency_counter_01),
	.read_latency_shift_reg_0(read_latency_shift_reg_02),
	.cp_ready(\seg_s1_agent|cp_ready~0_combout ),
	.WideOr1(\cmd_mux_005|WideOr1~combout ),
	.src_data_56(\cmd_mux_005|src_data[56]~combout ),
	.uav_write(uav_write),
	.av_readdata_pre_0(\seg_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(av_readdata_pre_13),
	.av_readdata_pre_4(av_readdata_pre_4),
	.av_readdata_pre_3(av_readdata_pre_33),
	.av_readdata_pre_2(av_readdata_pre_28),
	.av_readdata_pre_5(av_readdata_pre_5),
	.av_readdata_pre_7(av_readdata_pre_72),
	.av_readdata_pre_6(av_readdata_pre_62),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_71,readdata_61,readdata_5,readdata_4,readdata_32,readdata_21,readdata_12,readdata_01}),
	.clk(clk_clk));

processor_altera_merlin_slave_translator_4 seg_en_s1_translator(
	.reset(r_sync_rst),
	.rst1(rst1),
	.saved_grant_0(saved_grant_02),
	.src_valid(src_valid4),
	.src_valid1(src_valid5),
	.mem_used_1(mem_used_12),
	.always0(always02),
	.wait_latency_counter_1(wait_latency_counter_12),
	.wait_latency_counter_0(wait_latency_counter_02),
	.read_latency_shift_reg_0(\seg_en_s1_translator|read_latency_shift_reg[0]~q ),
	.cp_ready(\seg_en_s1_agent|cp_ready~0_combout ),
	.uav_write(uav_write),
	.WideOr1(\cmd_mux_004|WideOr1~combout ),
	.src_data_56(\cmd_mux_004|src_data[56]~combout ),
	.av_readdata_pre_0(\seg_en_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(av_readdata_pre_15),
	.av_readdata_pre_2(av_readdata_pre_29),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_27,readdata_14,readdata_02}),
	.clk(clk_clk));

processor_altera_merlin_slave_translator_1 led_s1_translator(
	.reset(r_sync_rst),
	.src_payload(src_payload),
	.rst1(rst1),
	.mem_used_1(mem_used_1),
	.always0(always0),
	.wait_latency_counter_1(wait_latency_counter_1),
	.wait_latency_counter_0(wait_latency_counter_0),
	.cp_ready(\led_s1_agent|cp_ready~0_combout ),
	.read_latency_shift_reg_0(\led_s1_translator|read_latency_shift_reg[0]~q ),
	.WideOr1(\cmd_mux_003|WideOr1~combout ),
	.src_data_56(\cmd_mux_003|src_data[56]~combout ),
	.read_latency_shift_reg(\led_s1_translator|read_latency_shift_reg~0_combout ),
	.av_readdata_pre_0(\led_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(av_readdata_pre_14),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_13,readdata_04}),
	.clk(clk_clk));

processor_altera_merlin_slave_translator_3 onchip_memory2_0_s1_translator(
	.reset(r_sync_rst),
	.rst1(rst1),
	.read_latency_shift_reg_0(read_latency_shift_reg_01),
	.mem_used_1(mem_used_13),
	.WideOr1(WideOr18),
	.mem(\onchip_memory2_0_s1_agent_rsp_fifo|mem~0_combout ),
	.read_latency_shift_reg(\onchip_memory2_0_s1_translator|read_latency_shift_reg~0_combout ),
	.clk(clk_clk));

processor_altera_merlin_slave_translator_2 nios2_gen2_0_debug_mem_slave_translator(
	.av_readdata({readdata_311,readdata_30,readdata_29,readdata_281,readdata_271,readdata_26,readdata_25,readdata_24,readdata_23,readdata_22,readdata_211,readdata_20,readdata_19,readdata_18,readdata_17,readdata_16,readdata_15,readdata_141,readdata_131,readdata_121,readdata_111,readdata_10,
readdata_9,readdata_8,readdata_7,readdata_6,readdata_52,readdata_42,readdata_3,readdata_2,readdata_1,readdata_0}),
	.reset(r_sync_rst),
	.rst1(rst1),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.write(\nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|write~0_combout ),
	.WideOr1(WideOr17),
	.mem(\nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|mem~0_combout ),
	.av_readdata_pre_0(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_22(av_readdata_pre_221),
	.av_readdata_pre_23(av_readdata_pre_23),
	.av_readdata_pre_24(av_readdata_pre_24),
	.av_readdata_pre_25(av_readdata_pre_25),
	.av_readdata_pre_26(av_readdata_pre_26),
	.av_readdata_pre_1(av_readdata_pre_11),
	.av_readdata_pre_4(av_readdata_pre_42),
	.av_readdata_pre_3(av_readdata_pre_31),
	.av_readdata_pre_2(av_readdata_pre_2),
	.av_readdata_pre_5(av_readdata_pre_52),
	.av_readdata_pre_14(av_readdata_pre_141),
	.av_readdata_pre_15(av_readdata_pre_151),
	.av_readdata_pre_11(av_readdata_pre_111),
	.av_readdata_pre_13(av_readdata_pre_131),
	.av_readdata_pre_16(av_readdata_pre_161),
	.av_readdata_pre_12(av_readdata_pre_121),
	.av_readdata_pre_10(av_readdata_pre_10),
	.av_readdata_pre_9(av_readdata_pre_9),
	.av_readdata_pre_8(av_readdata_pre_8),
	.av_readdata_pre_7(av_readdata_pre_7),
	.av_readdata_pre_6(av_readdata_pre_6),
	.av_readdata_pre_21(av_readdata_pre_211),
	.av_readdata_pre_20(av_readdata_pre_201),
	.av_readdata_pre_19(av_readdata_pre_191),
	.av_readdata_pre_18(av_readdata_pre_181),
	.av_readdata_pre_17(av_readdata_pre_171),
	.av_readdata_pre_27(av_readdata_pre_271),
	.av_readdata_pre_28(av_readdata_pre_281),
	.av_readdata_pre_29(av_readdata_pre_291),
	.av_readdata_pre_30(av_readdata_pre_30),
	.av_readdata_pre_31(av_readdata_pre_311),
	.clk(clk_clk));

processor_altera_merlin_slave_translator jtag_uart_0_avalon_jtag_slave_translator(
	.av_readdata_pre_22(av_readdata_pre_22),
	.av_readdata_pre_16(av_readdata_pre_16),
	.av_readdata_pre_21(av_readdata_pre_21),
	.av_readdata_pre_20(av_readdata_pre_20),
	.av_readdata_pre_19(av_readdata_pre_19),
	.av_readdata_pre_18(av_readdata_pre_18),
	.av_readdata_pre_17(av_readdata_pre_17),
	.reset(r_sync_rst),
	.rst1(rst1),
	.read_latency_shift_reg_0(\jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ),
	.sink_ready(\cmd_demux|sink_ready~4_combout ),
	.src_data_56(src_data_56),
	.WideOr1(WideOr16),
	.av_readdata_pre_0(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(av_readdata_pre_1),
	.av_readdata_pre_4(av_readdata_pre_43),
	.av_readdata_pre_3(av_readdata_pre_3),
	.av_readdata_pre_2(av_readdata_pre_27),
	.av_readdata_pre_5(av_readdata_pre_53),
	.av_readdata_pre_14(av_readdata_pre_142),
	.av_readdata_pre_15(av_readdata_pre_152),
	.av_readdata_pre_13(av_readdata_pre_132),
	.av_readdata_pre_12(av_readdata_pre_122),
	.av_readdata_pre_10(av_readdata_pre_101),
	.av_readdata_pre_9(av_readdata_pre_91),
	.av_readdata_pre_8(av_readdata_pre_81),
	.av_readdata_pre_7(av_readdata_pre_71),
	.av_readdata_pre_6(av_readdata_pre_61),
	.b_full(b_full),
	.read_0(read_0),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,rvalid,woverflow,gnd,b_non_empty,gnd,ac,av_readdata_9,av_readdata_8,av_readdata_7,av_readdata_6,av_readdata_5,av_readdata_4,av_readdata_3,av_readdata_2,av_readdata_1,av_readdata_0}),
	.b_full1(b_full1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_01(counter_reg_bit_01),
	.counter_reg_bit_51(counter_reg_bit_51),
	.counter_reg_bit_41(counter_reg_bit_41),
	.counter_reg_bit_31(counter_reg_bit_31),
	.counter_reg_bit_21(counter_reg_bit_21),
	.counter_reg_bit_11(counter_reg_bit_11),
	.clk(clk_clk));

processor_altera_merlin_master_translator nios2_gen2_0_data_master_translator(
	.reset(r_sync_rst),
	.d_write(d_write),
	.write_accepted1(\nios2_gen2_0_data_master_translator|write_accepted~q ),
	.rst1(rst1),
	.read_accepted1(\nios2_gen2_0_data_master_translator|read_accepted~q ),
	.d_read(d_read),
	.cp_valid(\nios2_gen2_0_data_master_agent|cp_valid~0_combout ),
	.WideOr1(WideOr12),
	.WideOr0(\cmd_demux|WideOr0~2_combout ),
	.av_waitrequest(nios2_gen2_0_data_master_waitrequest),
	.uav_read1(\nios2_gen2_0_data_master_translator|uav_read~combout ),
	.uav_write(uav_write),
	.clk(clk_clk));

processor_altera_merlin_master_translator_1 nios2_gen2_0_instruction_master_translator(
	.reset(r_sync_rst),
	.saved_grant_1(saved_grant_1),
	.rst1(rst1),
	.i_read(i_read),
	.read_accepted1(\nios2_gen2_0_instruction_master_translator|read_accepted~q ),
	.Equal4(\router_001|Equal4~0_combout ),
	.mem_used_1(mem_used_1),
	.saved_grant_11(saved_grant_11),
	.mem_used_11(mem_used_11),
	.saved_grant_12(saved_grant_12),
	.uav_read1(\nios2_gen2_0_instruction_master_translator|uav_read~combout ),
	.Equal6(\router_001|Equal6~1_combout ),
	.cp_ready(\led_s1_agent|cp_ready~0_combout ),
	.mem_used_12(mem_used_13),
	.mem_used_13(mem_used_14),
	.uav_waitrequest(\uart_0_s1_translator|uav_waitrequest~0_combout ),
	.sink_ready(\cmd_demux|sink_ready~4_combout ),
	.cp_ready1(\seg_s1_agent|cp_ready~0_combout ),
	.saved_grant_13(saved_grant_13),
	.WideOr1(WideOr13),
	.WideOr11(WideOr14),
	.Equal7(\router_001|Equal7~0_combout ),
	.saved_grant_14(\cmd_mux|saved_grant[1]~q ),
	.saved_grant_15(\cmd_mux_001|saved_grant[1]~q ),
	.write(\nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|write~0_combout ),
	.Equal1(\router_001|Equal1~1_combout ),
	.saved_grant_16(\cmd_mux_002|saved_grant[1]~q ),
	.Equal2(\router_001|Equal2~2_combout ),
	.src_channel_2(\router_001|src_channel[2]~2_combout ),
	.saved_grant_17(\cmd_mux_007|saved_grant[1]~q ),
	.Equal5(\router_001|Equal5~1_combout ),
	.cp_ready2(\seg_en_s1_agent|cp_ready~2_combout ),
	.Equal41(\router_001|Equal4~3_combout ),
	.always1(\router_001|always1~1_combout ),
	.cp_ready3(\sw_s1_agent|cp_ready~combout ),
	.clk(clk_clk));

processor_processor_mm_interconnect_0_cmd_mux cmd_mux(
	.W_alu_result_2(W_alu_result_2),
	.d_writedata_0(d_writedata_0),
	.r_sync_rst(r_sync_rst),
	.rst1(rst1),
	.Equal4(\router|Equal4~0_combout ),
	.cp_valid(\nios2_gen2_0_data_master_agent|cp_valid~0_combout ),
	.F_pc_0(F_pc_0),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.uav_read(\nios2_gen2_0_instruction_master_translator|uav_read~combout ),
	.Equal7(\router|Equal7~0_combout ),
	.sink_ready(\cmd_demux|sink_ready~4_combout ),
	.saved_grant_0(saved_grant_04),
	.saved_grant_1(\cmd_mux|saved_grant[1]~q ),
	.uav_read1(\nios2_gen2_0_data_master_translator|uav_read~combout ),
	.src_data_56(src_data_56),
	.src0_valid(\cmd_demux_001|src0_valid~0_combout ),
	.WideOr11(WideOr16),
	.src_data_38(src_data_382),
	.src_payload(src_payload50),
	.src_payload1(src_payload53),
	.src_payload2(src_payload54),
	.src_payload3(src_payload94),
	.src_payload4(src_payload100),
	.src_payload5(src_payload101),
	.src_payload6(src_payload102),
	.src_payload7(src_payload103),
	.clk_clk(clk_clk));

processor_processor_mm_interconnect_0_cmd_demux_1 cmd_demux_001(
	.rst1(rst1),
	.i_read(i_read),
	.read_accepted(\nios2_gen2_0_instruction_master_translator|read_accepted~q ),
	.cp_valid(\nios2_gen2_0_instruction_master_agent|cp_valid~combout ),
	.Equal1(\router_001|Equal1~0_combout ),
	.F_pc_10(F_pc_10),
	.F_pc_9(F_pc_9),
	.Equal4(\router_001|Equal4~0_combout ),
	.F_pc_2(F_pc_2),
	.Equal41(\router_001|Equal4~2_combout ),
	.uav_read(\nios2_gen2_0_instruction_master_translator|uav_read~combout ),
	.Equal6(\router_001|Equal6~1_combout ),
	.Equal7(\router_001|Equal7~0_combout ),
	.src_channel_2(\router_001|src_channel[2]~0_combout ),
	.Equal2(\router_001|Equal2~2_combout ),
	.src_channel_21(\router_001|src_channel[2]~1_combout ),
	.Equal5(\router_001|Equal5~1_combout ),
	.always1(\router_001|always1~1_combout ),
	.src5_valid(\cmd_demux_001|src5_valid~0_combout ),
	.src0_valid(\cmd_demux_001|src0_valid~0_combout ),
	.src1_valid(\cmd_demux_001|src1_valid~0_combout ),
	.src2_valid(\cmd_demux_001|src2_valid~0_combout ),
	.src6_valid(\cmd_demux_001|src6_valid~0_combout ),
	.src3_valid(\cmd_demux_001|src3_valid~2_combout ),
	.src4_valid(\cmd_demux_001|src4_valid~2_combout ),
	.src7_valid(\cmd_demux_001|src7_valid~2_combout ));

processor_processor_mm_interconnect_0_cmd_demux cmd_demux(
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_6(W_alu_result_6),
	.saved_grant_0(saved_grant_0),
	.rst1(rst1),
	.Equal4(\router|Equal4~0_combout ),
	.mem_used_1(mem_used_1),
	.saved_grant_01(saved_grant_01),
	.mem_used_11(mem_used_11),
	.saved_grant_02(saved_grant_02),
	.mem_used_12(mem_used_12),
	.Equal6(\router|Equal6~1_combout ),
	.cp_valid(\nios2_gen2_0_data_master_agent|cp_valid~1_combout ),
	.cp_ready(\led_s1_agent|cp_ready~0_combout ),
	.Equal5(\router|Equal5~1_combout ),
	.cp_ready1(\seg_en_s1_agent|cp_ready~0_combout ),
	.Equal1(\router|Equal1~1_combout ),
	.Equal7(\router|Equal7~0_combout ),
	.Equal2(\router|Equal2~2_combout ),
	.saved_grant_03(saved_grant_03),
	.mem_used_13(mem_used_13),
	.always1(\router|always1~1_combout ),
	.saved_grant_04(\cmd_mux_007|saved_grant[0]~q ),
	.mem_used_14(mem_used_14),
	.uav_waitrequest(\uart_0_s1_translator|uav_waitrequest~0_combout ),
	.av_waitrequest(av_waitrequest),
	.mem_used_15(mem_used_15),
	.sink_ready(\cmd_demux|sink_ready~4_combout ),
	.saved_grant_05(saved_grant_04),
	.saved_grant_06(saved_grant_05),
	.waitrequest(waitrequest),
	.mem_used_16(mem_used_16),
	.Equal41(\router|Equal4~1_combout ),
	.cp_ready2(\seg_s1_agent|cp_ready~0_combout ),
	.saved_grant_07(saved_grant_06),
	.mem_used_17(\sw_s1_agent_rsp_fifo|mem_used[1]~q ),
	.cp_ready3(\sw_s1_agent|cp_ready~0_combout ),
	.WideOr0(\cmd_demux|WideOr0~2_combout ),
	.src2_valid(\cmd_demux|src2_valid~2_combout ));

processor_processor_mm_interconnect_0_rsp_mux_1 rsp_mux_001(
	.q_a_0(q_a_0),
	.q_a_11(q_a_11),
	.read_latency_shift_reg_0(\jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo|mem[0][56]~q ),
	.read_latency_shift_reg_01(read_latency_shift_reg_01),
	.mem_74_01(mem_74_01),
	.mem_56_01(mem_56_01),
	.read_latency_shift_reg_02(\led_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_74_02(\led_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_02(\led_s1_agent_rsp_fifo|mem[0][56]~q ),
	.read_latency_shift_reg_03(\seg_en_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_74_03(\seg_en_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_03(\seg_en_s1_agent_rsp_fifo|mem[0][56]~q ),
	.read_latency_shift_reg_04(\sw_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_74_04(\sw_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_04(\sw_s1_agent_rsp_fifo|mem[0][56]~q ),
	.src1_valid(src1_valid),
	.src1_valid1(src1_valid1),
	.src1_valid2(src1_valid2),
	.src1_valid3(src1_valid3),
	.WideOr1(WideOr13),
	.src1_valid4(src1_valid4),
	.src_payload(src_payload3),
	.src_payload1(src_payload4),
	.WideOr11(WideOr14),
	.av_readdata_pre_0(\seg_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_01(\seg_en_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_02(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_03(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_04(\uart_0_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_05(\led_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_06(\sw_s1_translator|av_readdata_pre[0]~q ),
	.src_data_0(src_data_01),
	.src_data_01(src_data_02),
	.src_data_02(src_data_03),
	.av_readdata_pre_3(av_readdata_pre_3),
	.src_payload2(src_payload6),
	.src_payload3(src_payload7));

processor_processor_mm_interconnect_0_rsp_mux rsp_mux(
	.q_a_0(q_a_0),
	.q_a_22(q_a_22),
	.av_readdata_pre_22(av_readdata_pre_22),
	.q_a_23(q_a_23),
	.q_a_14(q_a_14),
	.q_a_15(q_a_15),
	.q_a_11(q_a_11),
	.q_a_13(q_a_13),
	.q_a_16(q_a_16),
	.av_readdata_pre_16(av_readdata_pre_16),
	.q_a_12(q_a_12),
	.q_a_10(q_a_10),
	.q_a_9(q_a_9),
	.q_a_8(q_a_8),
	.q_a_21(q_a_21),
	.av_readdata_pre_21(av_readdata_pre_21),
	.q_a_20(q_a_20),
	.av_readdata_pre_20(av_readdata_pre_20),
	.q_a_19(q_a_19),
	.av_readdata_pre_19(av_readdata_pre_19),
	.q_a_18(q_a_18),
	.av_readdata_pre_18(av_readdata_pre_18),
	.q_a_17(q_a_17),
	.av_readdata_pre_17(av_readdata_pre_17),
	.src0_valid(src0_valid),
	.src0_valid1(src0_valid1),
	.read_latency_shift_reg_0(read_latency_shift_reg_01),
	.mem_74_0(mem_74_01),
	.mem_56_0(mem_56_01),
	.src0_valid2(src0_valid2),
	.src0_valid3(src0_valid3),
	.WideOr11(WideOr1),
	.src0_valid4(src0_valid4),
	.src0_valid5(src0_valid5),
	.src0_valid6(\rsp_demux_006|src0_valid~0_combout ),
	.src0_valid7(src0_valid6),
	.WideOr12(WideOr11),
	.WideOr13(WideOr12),
	.av_readdata_pre_0(\seg_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_01(\seg_en_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_02(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_03(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_04(\uart_0_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_05(\led_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_06(\sw_s1_translator|av_readdata_pre[0]~q ),
	.src_data_0(src_data_0),
	.av_readdata_pre_221(av_readdata_pre_221),
	.av_readdata_pre_23(av_readdata_pre_23),
	.av_readdata_pre_14(av_readdata_pre_141),
	.av_readdata_pre_141(av_readdata_pre_142),
	.av_readdata_pre_15(av_readdata_pre_151),
	.av_readdata_pre_151(av_readdata_pre_152),
	.av_readdata_pre_11(av_readdata_pre_111),
	.av_readdata_pre_13(av_readdata_pre_131),
	.av_readdata_pre_131(av_readdata_pre_132),
	.av_readdata_pre_161(av_readdata_pre_161),
	.av_readdata_pre_12(av_readdata_pre_121),
	.av_readdata_pre_121(av_readdata_pre_122),
	.av_readdata_pre_10(av_readdata_pre_10),
	.av_readdata_pre_101(av_readdata_pre_101),
	.av_readdata_pre_9(av_readdata_pre_9),
	.av_readdata_pre_91(av_readdata_pre_91),
	.av_readdata_pre_92(av_readdata_pre_92),
	.av_readdata_pre_8(av_readdata_pre_8),
	.av_readdata_pre_81(av_readdata_pre_81),
	.av_readdata_pre_82(av_readdata_pre_82),
	.av_readdata_pre_211(av_readdata_pre_211),
	.av_readdata_pre_201(av_readdata_pre_201),
	.av_readdata_pre_191(av_readdata_pre_191),
	.av_readdata_pre_181(av_readdata_pre_181),
	.av_readdata_pre_171(av_readdata_pre_171),
	.src_data_8(src_data_8),
	.src_payload(src_payload38),
	.src_payload1(src_payload41),
	.src_payload2(src_payload43),
	.src_payload3(src_payload45),
	.src_payload4(src_payload47),
	.src_payload5(src_payload48),
	.src_payload6(src_payload49),
	.src_data_9(src_data_9),
	.src_payload7(src_payload60),
	.src_payload8(src_payload61),
	.src_payload9(src_payload62),
	.src_payload10(src_payload63),
	.src_payload11(src_payload64),
	.src_payload12(src_payload65),
	.src_payload13(src_payload66));

processor_processor_mm_interconnect_0_rsp_demux_7 rsp_demux_007(
	.read_latency_shift_reg_0(\uart_0_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\uart_0_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\uart_0_s1_agent_rsp_fifo|mem[0][56]~q ),
	.src0_valid(src0_valid6),
	.src1_valid(src1_valid4));

processor_processor_mm_interconnect_0_rsp_demux_6 rsp_demux_006(
	.read_latency_shift_reg_0(\sw_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\sw_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\sw_s1_agent_rsp_fifo|mem[0][56]~q ),
	.src0_valid(\rsp_demux_006|src0_valid~0_combout ));

processor_processor_mm_interconnect_0_rsp_demux_5 rsp_demux_005(
	.read_latency_shift_reg_0(read_latency_shift_reg_02),
	.mem_74_0(mem_74_02),
	.mem_56_0(mem_56_02),
	.src0_valid(src0_valid5),
	.src1_valid(src1_valid3));

processor_processor_mm_interconnect_0_rsp_demux_4 rsp_demux_004(
	.read_latency_shift_reg_0(\seg_en_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\seg_en_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\seg_en_s1_agent_rsp_fifo|mem[0][56]~q ),
	.src0_valid(src0_valid4));

processor_processor_mm_interconnect_0_rsp_demux_3 rsp_demux_003(
	.read_latency_shift_reg_0(\led_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\led_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\led_s1_agent_rsp_fifo|mem[0][56]~q ),
	.src0_valid(src0_valid3));

processor_processor_mm_interconnect_0_rsp_demux_2 rsp_demux_002(
	.read_latency_shift_reg_0(read_latency_shift_reg_01),
	.mem_74_0(mem_74_01),
	.mem_56_0(mem_56_01),
	.src0_valid(src0_valid2),
	.src1_valid(src1_valid2));

processor_processor_mm_interconnect_0_rsp_demux_1 rsp_demux_001(
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.mem_74_0(mem_74_0),
	.mem_56_0(mem_56_0),
	.src0_valid(src0_valid1),
	.src1_valid(src1_valid1));

processor_processor_mm_interconnect_0_rsp_demux rsp_demux(
	.read_latency_shift_reg_0(\jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo|mem[0][56]~q ),
	.src0_valid(src0_valid),
	.src1_valid(src1_valid));

processor_processor_mm_interconnect_0_cmd_mux_7 cmd_mux_007(
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_2(W_alu_result_2),
	.W_alu_result_3(W_alu_result_3),
	.d_writedata_0(d_writedata_0),
	.r_sync_rst(r_sync_rst),
	.rst1(rst1),
	.F_pc_2(F_pc_2),
	.cp_valid(\nios2_gen2_0_data_master_agent|cp_valid~0_combout ),
	.F_pc_1(F_pc_1),
	.F_pc_0(F_pc_0),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.uav_read(\nios2_gen2_0_instruction_master_translator|uav_read~combout ),
	.Equal2(\router|Equal2~2_combout ),
	.saved_grant_0(\cmd_mux_007|saved_grant[0]~q ),
	.mem_used_1(mem_used_14),
	.uav_waitrequest(\uart_0_s1_translator|uav_waitrequest~0_combout ),
	.saved_grant_1(\cmd_mux_007|saved_grant[1]~q ),
	.uav_read1(\nios2_gen2_0_data_master_translator|uav_read~combout ),
	.d_writedata_9(d_writedata_9),
	.src_payload(src_payload5),
	.src_data_38(src_data_38),
	.src_data_39(src_data_39),
	.src_data_40(src_data_40),
	.WideOr11(WideOr15),
	.src_data_56(src_data_561),
	.src_payload1(src_payload8),
	.src_payload2(src_payload9),
	.src_payload3(src_payload10),
	.src_payload4(src_payload11),
	.src_payload5(src_payload12),
	.src_payload6(src_payload13),
	.src_payload7(src_payload14),
	.src_payload8(src_payload15),
	.d_writedata_8(d_writedata_8),
	.src_payload9(src_payload68),
	.src7_valid(\cmd_demux_001|src7_valid~2_combout ),
	.clk_clk(clk_clk));

processor_processor_mm_interconnect_0_cmd_mux_6 cmd_mux_006(
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_6(W_alu_result_6),
	.r_sync_rst(r_sync_rst),
	.rst1(rst1),
	.cp_valid(\nios2_gen2_0_instruction_master_agent|cp_valid~combout ),
	.Equal4(\router|Equal4~0_combout ),
	.cp_valid1(\nios2_gen2_0_data_master_agent|cp_valid~0_combout ),
	.Equal41(\router_001|Equal4~2_combout ),
	.uav_read(\nios2_gen2_0_instruction_master_translator|uav_read~combout ),
	.always1(\router|always1~0_combout ),
	.always11(\router|always1~1_combout ),
	.saved_grant_0(saved_grant_06),
	.always12(\router_001|always1~0_combout ),
	.saved_grant_1(saved_grant_13),
	.src_valid(\cmd_mux_006|src_valid~2_combout ),
	.src_valid1(\cmd_mux_006|src_valid~4_combout ),
	.always13(\router_001|always1~1_combout ),
	.cp_ready(\sw_s1_agent|cp_ready~combout ),
	.uav_read1(\nios2_gen2_0_data_master_translator|uav_read~combout ),
	.WideOr11(\cmd_mux_006|WideOr1~combout ),
	.src_data_56(\cmd_mux_006|src_data[56]~combout ),
	.src6_valid(\cmd_demux_001|src6_valid~0_combout ),
	.clk_clk(clk_clk));

processor_processor_mm_interconnect_0_cmd_mux_5 cmd_mux_005(
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_6(W_alu_result_6),
	.r_sync_rst(r_sync_rst),
	.d_write(d_write),
	.write_accepted(\nios2_gen2_0_data_master_translator|write_accepted~q ),
	.rst1(rst1),
	.cp_valid(\nios2_gen2_0_instruction_master_agent|cp_valid~combout ),
	.F_pc_2(F_pc_2),
	.Equal4(\router|Equal4~0_combout ),
	.cp_valid1(\nios2_gen2_0_data_master_agent|cp_valid~0_combout ),
	.saved_grant_0(saved_grant_01),
	.src_payload(src_payload1),
	.saved_grant_1(saved_grant_11),
	.Equal41(\router_001|Equal4~2_combout ),
	.src_valid(src_valid2),
	.src_valid1(src_valid3),
	.uav_read(\nios2_gen2_0_instruction_master_translator|uav_read~combout ),
	.Equal42(\router|Equal4~1_combout ),
	.uav_read1(\nios2_gen2_0_data_master_translator|uav_read~combout ),
	.src5_valid(\cmd_demux_001|src5_valid~0_combout ),
	.write(\seg_s1_agent_rsp_fifo|write~1_combout ),
	.WideOr11(\cmd_mux_005|WideOr1~combout ),
	.src_data_56(\cmd_mux_005|src_data[56]~combout ),
	.clk_clk(clk_clk));

processor_processor_mm_interconnect_0_cmd_mux_4 cmd_mux_004(
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_6(W_alu_result_6),
	.r_sync_rst(r_sync_rst),
	.d_write(d_write),
	.write_accepted(\nios2_gen2_0_data_master_translator|write_accepted~q ),
	.rst1(rst1),
	.cp_valid(\nios2_gen2_0_instruction_master_agent|cp_valid~combout ),
	.Equal4(\router_001|Equal4~0_combout ),
	.F_pc_2(F_pc_2),
	.F_pc_3(F_pc_3),
	.F_pc_4(F_pc_4),
	.Equal41(\router|Equal4~0_combout ),
	.cp_valid1(\nios2_gen2_0_data_master_agent|cp_valid~0_combout ),
	.saved_grant_0(saved_grant_02),
	.src_payload(src_payload2),
	.saved_grant_1(saved_grant_12),
	.src_valid(src_valid4),
	.src_valid1(src_valid5),
	.uav_read(\nios2_gen2_0_instruction_master_translator|uav_read~combout ),
	.Equal5(\router|Equal5~1_combout ),
	.cp_ready(\seg_en_s1_agent|cp_ready~2_combout ),
	.uav_read1(\nios2_gen2_0_data_master_translator|uav_read~combout ),
	.WideOr11(\cmd_mux_004|WideOr1~combout ),
	.src_data_56(\cmd_mux_004|src_data[56]~combout ),
	.src_valid2(\cmd_mux_004|src_valid~6_combout ),
	.src4_valid(\cmd_demux_001|src4_valid~2_combout ),
	.clk_clk(clk_clk));

processor_processor_mm_interconnect_0_cmd_mux_3 cmd_mux_003(
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_6(W_alu_result_6),
	.r_sync_rst(r_sync_rst),
	.saved_grant_0(saved_grant_0),
	.d_write(d_write),
	.write_accepted(\nios2_gen2_0_data_master_translator|write_accepted~q ),
	.src_payload(src_payload),
	.saved_grant_1(saved_grant_1),
	.rst1(rst1),
	.cp_valid(\nios2_gen2_0_instruction_master_agent|cp_valid~combout ),
	.Equal4(\router_001|Equal4~0_combout ),
	.F_pc_2(F_pc_2),
	.F_pc_3(F_pc_3),
	.F_pc_4(F_pc_4),
	.src_valid(src_valid),
	.Equal41(\router|Equal4~0_combout ),
	.cp_valid1(\nios2_gen2_0_data_master_agent|cp_valid~0_combout ),
	.src_valid1(src_valid1),
	.mem_used_1(mem_used_1),
	.Equal6(\router|Equal6~1_combout ),
	.uav_read(\nios2_gen2_0_instruction_master_translator|uav_read~combout ),
	.cp_ready(\led_s1_agent|cp_ready~0_combout ),
	.WideOr11(\cmd_mux_003|WideOr1~combout ),
	.uav_read1(\nios2_gen2_0_data_master_translator|uav_read~combout ),
	.src_data_56(\cmd_mux_003|src_data[56]~combout ),
	.src3_valid(\cmd_demux_001|src3_valid~2_combout ),
	.clk_clk(clk_clk));

processor_processor_mm_interconnect_0_cmd_mux_2 cmd_mux_002(
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_14(W_alu_result_14),
	.W_alu_result_13(W_alu_result_13),
	.W_alu_result_12(W_alu_result_12),
	.W_alu_result_11(W_alu_result_11),
	.W_alu_result_10(W_alu_result_10),
	.W_alu_result_9(W_alu_result_9),
	.W_alu_result_8(W_alu_result_8),
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_6(W_alu_result_6),
	.W_alu_result_2(W_alu_result_2),
	.W_alu_result_3(W_alu_result_3),
	.d_writedata_24(d_writedata_24),
	.d_writedata_25(d_writedata_25),
	.d_writedata_26(d_writedata_26),
	.d_writedata_27(d_writedata_27),
	.d_writedata_28(d_writedata_28),
	.d_writedata_29(d_writedata_29),
	.d_writedata_30(d_writedata_30),
	.d_writedata_31(d_writedata_31),
	.d_writedata_0(d_writedata_0),
	.r_sync_rst(r_sync_rst),
	.rst1(rst1),
	.F_pc_5(F_pc_5),
	.F_pc_12(F_pc_12),
	.F_pc_11(F_pc_11),
	.F_pc_10(F_pc_10),
	.F_pc_9(F_pc_9),
	.F_pc_8(F_pc_8),
	.F_pc_7(F_pc_7),
	.F_pc_6(F_pc_6),
	.F_pc_2(F_pc_2),
	.F_pc_3(F_pc_3),
	.F_pc_4(F_pc_4),
	.F_pc_1(F_pc_1),
	.F_pc_0(F_pc_0),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.saved_grant_0(saved_grant_03),
	.mem_used_1(mem_used_13),
	.saved_grant_1(\cmd_mux_002|saved_grant[1]~q ),
	.d_writedata_9(d_writedata_9),
	.src2_valid(\cmd_demux|src2_valid~2_combout ),
	.src2_valid1(\cmd_demux_001|src2_valid~0_combout ),
	.WideOr11(WideOr18),
	.src_payload(src_payload16),
	.src_data_38(src_data_381),
	.src_data_39(src_data_391),
	.src_data_40(src_data_401),
	.src_data_41(src_data_41),
	.src_data_42(src_data_42),
	.src_data_43(src_data_43),
	.src_data_44(src_data_44),
	.src_data_45(src_data_45),
	.src_data_46(src_data_461),
	.src_data_47(src_data_47),
	.src_data_48(src_data_48),
	.src_data_49(src_data_49),
	.src_data_50(src_data_50),
	.d_byteenable_0(d_byteenable_0),
	.src_data_32(src_data_32),
	.d_writedata_22(d_writedata_22),
	.src_payload1(src_payload17),
	.d_byteenable_2(d_byteenable_2),
	.src_data_34(src_data_34),
	.d_writedata_23(d_writedata_23),
	.src_payload2(src_payload18),
	.src_payload3(src_payload19),
	.d_byteenable_3(d_byteenable_3),
	.src_data_35(src_data_35),
	.src_payload4(src_payload20),
	.src_payload5(src_payload21),
	.src_payload6(src_payload22),
	.src_payload7(src_payload23),
	.src_payload8(src_payload24),
	.src_payload9(src_payload25),
	.src_payload10(src_payload26),
	.d_writedata_14(d_writedata_14),
	.src_payload11(src_payload27),
	.d_byteenable_1(d_byteenable_1),
	.src_data_33(src_data_33),
	.d_writedata_15(d_writedata_15),
	.src_payload12(src_payload28),
	.d_writedata_11(d_writedata_11),
	.src_payload13(src_payload29),
	.d_writedata_13(d_writedata_13),
	.src_payload14(src_payload30),
	.d_writedata_16(d_writedata_16),
	.src_payload15(src_payload31),
	.d_writedata_12(d_writedata_12),
	.src_payload16(src_payload32),
	.d_writedata_10(d_writedata_10),
	.src_payload17(src_payload33),
	.src_payload18(src_payload34),
	.d_writedata_8(d_writedata_8),
	.src_payload19(src_payload35),
	.src_payload20(src_payload36),
	.src_payload21(src_payload37),
	.d_writedata_21(d_writedata_21),
	.src_payload22(src_payload39),
	.d_writedata_20(d_writedata_20),
	.src_payload23(src_payload40),
	.d_writedata_19(d_writedata_19),
	.src_payload24(src_payload42),
	.d_writedata_18(d_writedata_18),
	.src_payload25(src_payload44),
	.d_writedata_17(d_writedata_17),
	.src_payload26(src_payload46),
	.src_payload27(src_payload55),
	.src_payload28(src_payload56),
	.src_payload29(src_payload57),
	.src_payload30(src_payload58),
	.src_payload31(src_payload59),
	.clk_clk(clk_clk));

processor_processor_mm_interconnect_0_cmd_mux_1 cmd_mux_001(
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_10(W_alu_result_10),
	.W_alu_result_9(W_alu_result_9),
	.W_alu_result_8(W_alu_result_8),
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_6(W_alu_result_6),
	.W_alu_result_2(W_alu_result_2),
	.W_alu_result_3(W_alu_result_3),
	.d_writedata_24(d_writedata_24),
	.d_writedata_25(d_writedata_25),
	.d_writedata_26(d_writedata_26),
	.d_writedata_27(d_writedata_27),
	.d_writedata_28(d_writedata_28),
	.d_writedata_29(d_writedata_29),
	.d_writedata_30(d_writedata_30),
	.d_writedata_31(d_writedata_31),
	.d_writedata_0(d_writedata_0),
	.r_sync_rst(r_sync_rst),
	.rst1(rst1),
	.F_pc_5(F_pc_5),
	.F_pc_8(F_pc_8),
	.F_pc_7(F_pc_7),
	.F_pc_6(F_pc_6),
	.F_pc_2(F_pc_2),
	.F_pc_3(F_pc_3),
	.F_pc_4(F_pc_4),
	.cp_valid(\nios2_gen2_0_data_master_agent|cp_valid~0_combout ),
	.F_pc_1(F_pc_1),
	.F_pc_0(F_pc_0),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.Equal1(\router|Equal1~1_combout ),
	.saved_grant_0(saved_grant_05),
	.waitrequest(waitrequest),
	.mem_used_1(mem_used_16),
	.saved_grant_1(\cmd_mux_001|saved_grant[1]~q ),
	.d_writedata_9(d_writedata_9),
	.src1_valid(\cmd_demux_001|src1_valid~0_combout ),
	.WideOr11(WideOr17),
	.hbreak_enabled(hbreak_enabled),
	.src_data_46(src_data_46),
	.d_byteenable_0(d_byteenable_0),
	.d_writedata_22(d_writedata_22),
	.d_byteenable_2(d_byteenable_2),
	.d_writedata_23(d_writedata_23),
	.d_byteenable_3(d_byteenable_3),
	.d_writedata_14(d_writedata_14),
	.d_byteenable_1(d_byteenable_1),
	.d_writedata_15(d_writedata_15),
	.d_writedata_11(d_writedata_11),
	.d_writedata_13(d_writedata_13),
	.d_writedata_16(d_writedata_16),
	.d_writedata_12(d_writedata_12),
	.d_writedata_10(d_writedata_10),
	.d_writedata_8(d_writedata_8),
	.d_writedata_21(d_writedata_21),
	.d_writedata_20(d_writedata_20),
	.d_writedata_19(d_writedata_19),
	.d_writedata_18(d_writedata_18),
	.d_writedata_17(d_writedata_17),
	.src_payload(src_payload51),
	.src_payload1(src_payload52),
	.src_data_38(src_data_383),
	.src_data_39(src_data_392),
	.src_data_40(src_data_402),
	.src_data_41(src_data_411),
	.src_data_42(src_data_421),
	.src_data_43(src_data_431),
	.src_data_44(src_data_441),
	.src_data_45(src_data_451),
	.src_data_32(src_data_321),
	.src_payload2(src_payload67),
	.src_payload3(src_payload69),
	.src_payload4(src_payload70),
	.src_payload5(src_payload71),
	.src_data_34(src_data_341),
	.src_payload6(src_payload72),
	.src_payload7(src_payload73),
	.src_data_35(src_data_351),
	.src_payload8(src_payload74),
	.src_payload9(src_payload75),
	.src_payload10(src_payload76),
	.src_payload11(src_payload77),
	.src_payload12(src_payload78),
	.src_data_33(src_data_331),
	.src_payload13(src_payload79),
	.src_payload14(src_payload80),
	.src_payload15(src_payload81),
	.src_payload16(src_payload82),
	.src_payload17(src_payload83),
	.src_payload18(src_payload84),
	.src_payload19(src_payload85),
	.src_payload20(src_payload86),
	.src_payload21(src_payload87),
	.src_payload22(src_payload88),
	.src_payload23(src_payload89),
	.src_payload24(src_payload90),
	.src_payload25(src_payload91),
	.src_payload26(src_payload92),
	.src_payload27(src_payload93),
	.src_payload28(src_payload95),
	.src_payload29(src_payload96),
	.src_payload30(src_payload97),
	.src_payload31(src_payload98),
	.src_payload32(src_payload99),
	.clk_clk(clk_clk));

endmodule

module processor_altera_avalon_sc_fifo (
	reset,
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	av_waitrequest,
	mem_used_1,
	sink_ready,
	saved_grant_1,
	src_data_56,
	WideOr1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	read_latency_shift_reg_0;
output 	mem_74_0;
output 	mem_56_0;
input 	av_waitrequest;
output 	mem_used_1;
input 	sink_ready;
input 	saved_grant_1;
input 	src_data_56;
input 	WideOr1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem[1][74]~q ;
wire \mem~0_combout ;
wire \mem_used[0]~3_combout ;
wire \mem_used[0]~4_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem[1][56]~q ;
wire \mem~1_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~2_combout ;


dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][56] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_56_0),
	.prn(vcc));
defparam \mem[0][56] .is_wysiwyg = "true";
defparam \mem[0][56] .power_up = "low";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclone10lp_lcell_comb \mem~0 (
	.dataa(\mem[1][74]~q ),
	.datab(saved_grant_1),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~0_combout ),
	.cout());
defparam \mem~0 .lut_mask = 16'hAACC;
defparam \mem~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_used[0]~3 (
	.dataa(\mem_used[0]~q ),
	.datab(mem_used_1),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hEEFF;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_used[0]~4 (
	.dataa(\mem_used[0]~3_combout ),
	.datab(sink_ready),
	.datac(src_data_56),
	.datad(WideOr1),
	.cin(gnd),
	.combout(\mem_used[0]~4_combout ),
	.cout());
defparam \mem_used[0]~4 .lut_mask = 16'hFFFE;
defparam \mem_used[0]~4 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclone10lp_lcell_comb \mem_used[1]~0 (
	.dataa(\mem_used[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hFF55;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

dffeas \mem[1][56] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][56]~q ),
	.prn(vcc));
defparam \mem[1][56] .is_wysiwyg = "true";
defparam \mem[1][56] .power_up = "low";

cyclone10lp_lcell_comb \mem~1 (
	.dataa(\mem[1][56]~q ),
	.datab(src_data_56),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~1_combout ),
	.cout());
defparam \mem~1 .lut_mask = 16'hAACC;
defparam \mem~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_used[1]~1 (
	.dataa(av_waitrequest),
	.datab(src_data_56),
	.datac(WideOr1),
	.datad(\mem_used[1]~0_combout ),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hFEFF;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_used[1]~2 (
	.dataa(\mem_used[1]~1_combout ),
	.datab(mem_used_1),
	.datac(read_latency_shift_reg_0),
	.datad(\mem_used[0]~q ),
	.cin(gnd),
	.combout(\mem_used[1]~2_combout ),
	.cout());
defparam \mem_used[1]~2 .lut_mask = 16'hEFFF;
defparam \mem_used[1]~2 .sum_lutc_input = "datac";

endmodule

module processor_altera_avalon_sc_fifo_1 (
	reset,
	saved_grant_1,
	mem_used_1,
	cp_ready,
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	WideOr1,
	src_data_56,
	read_latency_shift_reg,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	saved_grant_1;
output 	mem_used_1;
input 	cp_ready;
input 	read_latency_shift_reg_0;
output 	mem_74_0;
output 	mem_56_0;
input 	WideOr1;
input 	src_data_56;
input 	read_latency_shift_reg;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~3_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~2_combout ;
wire \mem[1][74]~q ;
wire \mem~0_combout ;
wire \mem[1][56]~q ;
wire \mem~1_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][56] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_56_0),
	.prn(vcc));
defparam \mem[0][56] .is_wysiwyg = "true";
defparam \mem[0][56] .power_up = "low";

cyclone10lp_lcell_comb \mem_used[0]~3 (
	.dataa(read_latency_shift_reg),
	.datab(\mem_used[0]~q ),
	.datac(mem_used_1),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hFEFF;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclone10lp_lcell_comb \mem_used[1]~0 (
	.dataa(\mem_used[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hFF55;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_used[1]~1 (
	.dataa(WideOr1),
	.datab(cp_ready),
	.datac(src_data_56),
	.datad(\mem_used[1]~0_combout ),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hFEFF;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_used[1]~2 (
	.dataa(\mem_used[1]~1_combout ),
	.datab(mem_used_1),
	.datac(read_latency_shift_reg_0),
	.datad(\mem_used[0]~q ),
	.cin(gnd),
	.combout(\mem_used[1]~2_combout ),
	.cout());
defparam \mem_used[1]~2 .lut_mask = 16'hEFFF;
defparam \mem_used[1]~2 .sum_lutc_input = "datac";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclone10lp_lcell_comb \mem~0 (
	.dataa(\mem[1][74]~q ),
	.datab(saved_grant_1),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~0_combout ),
	.cout());
defparam \mem~0 .lut_mask = 16'hAACC;
defparam \mem~0 .sum_lutc_input = "datac";

dffeas \mem[1][56] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][56]~q ),
	.prn(vcc));
defparam \mem[1][56] .is_wysiwyg = "true";
defparam \mem[1][56] .power_up = "low";

cyclone10lp_lcell_comb \mem~1 (
	.dataa(\mem[1][56]~q ),
	.datab(src_data_56),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~1_combout ),
	.cout());
defparam \mem~1 .lut_mask = 16'hAACC;
defparam \mem~1 .sum_lutc_input = "datac";

endmodule

module processor_altera_avalon_sc_fifo_2 (
	reset,
	uav_read,
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	saved_grant_0,
	waitrequest,
	mem_used_1,
	saved_grant_1,
	write,
	uav_read1,
	WideOr1,
	mem,
	rf_source_valid,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	uav_read;
input 	read_latency_shift_reg_0;
output 	mem_74_0;
output 	mem_56_0;
input 	saved_grant_0;
input 	waitrequest;
output 	mem_used_1;
input 	saved_grant_1;
output 	write;
input 	uav_read1;
input 	WideOr1;
output 	mem;
input 	rf_source_valid;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem[1][74]~q ;
wire \mem~1_combout ;
wire \mem_used[0]~3_combout ;
wire \mem_used[0]~4_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem[1][56]~q ;
wire \mem~2_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~2_combout ;


dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][56] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_56_0),
	.prn(vcc));
defparam \mem[0][56] .is_wysiwyg = "true";
defparam \mem[0][56] .power_up = "low";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclone10lp_lcell_comb \write~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(waitrequest),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(write),
	.cout());
defparam \write~0 .lut_mask = 16'h0FFF;
defparam \write~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem~0 (
	.dataa(uav_read),
	.datab(uav_read1),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(mem),
	.cout());
defparam \mem~0 .lut_mask = 16'hFFFE;
defparam \mem~0 .sum_lutc_input = "datac";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclone10lp_lcell_comb \mem~1 (
	.dataa(\mem[1][74]~q ),
	.datab(saved_grant_1),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~1_combout ),
	.cout());
defparam \mem~1 .lut_mask = 16'hAACC;
defparam \mem~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_used[0]~3 (
	.dataa(\mem_used[0]~q ),
	.datab(mem_used_1),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hEEFF;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_used[0]~4 (
	.dataa(\mem_used[0]~3_combout ),
	.datab(write),
	.datac(WideOr1),
	.datad(mem),
	.cin(gnd),
	.combout(\mem_used[0]~4_combout ),
	.cout());
defparam \mem_used[0]~4 .lut_mask = 16'hFFFE;
defparam \mem_used[0]~4 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclone10lp_lcell_comb \mem_used[1]~0 (
	.dataa(\mem_used[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hFF55;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

dffeas \mem[1][56] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][56]~q ),
	.prn(vcc));
defparam \mem[1][56] .is_wysiwyg = "true";
defparam \mem[1][56] .power_up = "low";

cyclone10lp_lcell_comb \mem~2 (
	.dataa(\mem[1][56]~q ),
	.datab(mem),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~2_combout ),
	.cout());
defparam \mem~2 .lut_mask = 16'hAACC;
defparam \mem~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_used[1]~1 (
	.dataa(mem_used_1),
	.datab(gnd),
	.datac(read_latency_shift_reg_0),
	.datad(\mem_used[0]~q ),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hAFFF;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_used[1]~2 (
	.dataa(\mem_used[1]~1_combout ),
	.datab(rf_source_valid),
	.datac(\mem_used[1]~0_combout ),
	.datad(waitrequest),
	.cin(gnd),
	.combout(\mem_used[1]~2_combout ),
	.cout());
defparam \mem_used[1]~2 .lut_mask = 16'hEFFF;
defparam \mem_used[1]~2 .sum_lutc_input = "datac";

endmodule

module processor_altera_avalon_sc_fifo_3 (
	reset,
	rst1,
	uav_read,
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	saved_grant_0,
	mem_used_1,
	saved_grant_1,
	uav_read1,
	WideOr1,
	mem,
	read_latency_shift_reg,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	rst1;
input 	uav_read;
input 	read_latency_shift_reg_0;
output 	mem_74_0;
output 	mem_56_0;
input 	saved_grant_0;
output 	mem_used_1;
input 	saved_grant_1;
input 	uav_read1;
input 	WideOr1;
output 	mem;
input 	read_latency_shift_reg;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem[1][74]~q ;
wire \mem~1_combout ;
wire \mem_used[0]~3_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem[1][56]~q ;
wire \mem~2_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~2_combout ;


dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][56] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_56_0),
	.prn(vcc));
defparam \mem[0][56] .is_wysiwyg = "true";
defparam \mem[0][56] .power_up = "low";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclone10lp_lcell_comb \mem~0 (
	.dataa(uav_read),
	.datab(uav_read1),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(mem),
	.cout());
defparam \mem~0 .lut_mask = 16'hFFFE;
defparam \mem~0 .sum_lutc_input = "datac";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclone10lp_lcell_comb \mem~1 (
	.dataa(\mem[1][74]~q ),
	.datab(saved_grant_1),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~1_combout ),
	.cout());
defparam \mem~1 .lut_mask = 16'hAACC;
defparam \mem~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_used[0]~3 (
	.dataa(read_latency_shift_reg),
	.datab(\mem_used[0]~q ),
	.datac(mem_used_1),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hFEFF;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclone10lp_lcell_comb \mem_used[1]~0 (
	.dataa(\mem_used[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hFF55;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

dffeas \mem[1][56] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][56]~q ),
	.prn(vcc));
defparam \mem[1][56] .is_wysiwyg = "true";
defparam \mem[1][56] .power_up = "low";

cyclone10lp_lcell_comb \mem~2 (
	.dataa(\mem[1][56]~q ),
	.datab(mem),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~2_combout ),
	.cout());
defparam \mem~2 .lut_mask = 16'hAACC;
defparam \mem~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_used[1]~1 (
	.dataa(rst1),
	.datab(WideOr1),
	.datac(mem),
	.datad(\mem_used[1]~0_combout ),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hFEFF;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_used[1]~2 (
	.dataa(\mem_used[1]~1_combout ),
	.datab(mem_used_1),
	.datac(read_latency_shift_reg_0),
	.datad(\mem_used[0]~q ),
	.cin(gnd),
	.combout(\mem_used[1]~2_combout ),
	.cout());
defparam \mem_used[1]~2 .lut_mask = 16'hEFFF;
defparam \mem_used[1]~2 .sum_lutc_input = "datac";

endmodule

module processor_altera_avalon_sc_fifo_4 (
	reset,
	saved_grant_0,
	saved_grant_1,
	src_valid,
	mem_used_1,
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	cp_ready,
	src_data_56,
	src_valid1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	saved_grant_0;
input 	saved_grant_1;
input 	src_valid;
output 	mem_used_1;
input 	read_latency_shift_reg_0;
output 	mem_74_0;
output 	mem_56_0;
input 	cp_ready;
input 	src_data_56;
input 	src_valid1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~3_combout ;
wire \write~0_combout ;
wire \mem_used[0]~4_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~2_combout ;
wire \mem[1][74]~q ;
wire \mem~0_combout ;
wire \mem[1][56]~q ;
wire \mem~1_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~1_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][56] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~1_combout ),
	.q(mem_56_0),
	.prn(vcc));
defparam \mem[0][56] .is_wysiwyg = "true";
defparam \mem[0][56] .power_up = "low";

cyclone10lp_lcell_comb \mem_used[0]~3 (
	.dataa(\mem_used[0]~q ),
	.datab(mem_used_1),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hEEFF;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \write~0 (
	.dataa(src_data_56),
	.datab(src_valid),
	.datac(saved_grant_0),
	.datad(src_valid1),
	.cin(gnd),
	.combout(\write~0_combout ),
	.cout());
defparam \write~0 .lut_mask = 16'hFFFE;
defparam \write~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_used[0]~4 (
	.dataa(\mem_used[0]~3_combout ),
	.datab(cp_ready),
	.datac(\write~0_combout ),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem_used[0]~4_combout ),
	.cout());
defparam \mem_used[0]~4 .lut_mask = 16'hFEFF;
defparam \mem_used[0]~4 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclone10lp_lcell_comb \mem_used[1]~0 (
	.dataa(mem_used_1),
	.datab(gnd),
	.datac(read_latency_shift_reg_0),
	.datad(\mem_used[0]~q ),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hAFFF;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_used[1]~1 (
	.dataa(\mem_used[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hFF55;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_used[1]~2 (
	.dataa(\mem_used[1]~0_combout ),
	.datab(cp_ready),
	.datac(\write~0_combout ),
	.datad(\mem_used[1]~1_combout ),
	.cin(gnd),
	.combout(\mem_used[1]~2_combout ),
	.cout());
defparam \mem_used[1]~2 .lut_mask = 16'hFEFF;
defparam \mem_used[1]~2 .sum_lutc_input = "datac";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclone10lp_lcell_comb \mem~0 (
	.dataa(\mem[1][74]~q ),
	.datab(saved_grant_1),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~0_combout ),
	.cout());
defparam \mem~0 .lut_mask = 16'hAACC;
defparam \mem~0 .sum_lutc_input = "datac";

dffeas \mem[1][56] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][56]~q ),
	.prn(vcc));
defparam \mem[1][56] .is_wysiwyg = "true";
defparam \mem[1][56] .power_up = "low";

cyclone10lp_lcell_comb \mem~1 (
	.dataa(\mem[1][56]~q ),
	.datab(src_data_56),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~1_combout ),
	.cout());
defparam \mem~1 .lut_mask = 16'hAACC;
defparam \mem~1 .sum_lutc_input = "datac";

endmodule

module processor_altera_avalon_sc_fifo_5 (
	reset,
	rst1,
	saved_grant_1,
	src_valid,
	src_valid1,
	mem_used_1,
	always0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	cp_ready,
	write,
	WideOr1,
	src_data_56,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	rst1;
input 	saved_grant_1;
input 	src_valid;
input 	src_valid1;
output 	mem_used_1;
input 	always0;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	read_latency_shift_reg_0;
output 	mem_74_0;
output 	mem_56_0;
input 	cp_ready;
output 	write;
input 	WideOr1;
input 	src_data_56;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~3_combout ;
wire \mem_used[0]~4_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~2_combout ;
wire \mem[1][74]~q ;
wire \mem~0_combout ;
wire \mem[1][56]~q ;
wire \mem~1_combout ;
wire \write~0_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][56] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_56_0),
	.prn(vcc));
defparam \mem[0][56] .is_wysiwyg = "true";
defparam \mem[0][56] .power_up = "low";

cyclone10lp_lcell_comb \write~1 (
	.dataa(mem_used_1),
	.datab(always0),
	.datac(wait_latency_counter_0),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(write),
	.cout());
defparam \write~1 .lut_mask = 16'hFF7D;
defparam \write~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_used[0]~3 (
	.dataa(\mem_used[0]~q ),
	.datab(mem_used_1),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hEEFF;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_used[0]~4 (
	.dataa(\mem_used[0]~3_combout ),
	.datab(src_data_56),
	.datac(write),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_used[0]~4_combout ),
	.cout());
defparam \mem_used[0]~4 .lut_mask = 16'hFEFE;
defparam \mem_used[0]~4 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclone10lp_lcell_comb \mem_used[1]~0 (
	.dataa(\mem_used[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hFF55;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_used[1]~1 (
	.dataa(WideOr1),
	.datab(cp_ready),
	.datac(\mem_used[1]~0_combout ),
	.datad(src_data_56),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hFFEF;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_used[1]~2 (
	.dataa(\mem_used[1]~1_combout ),
	.datab(mem_used_1),
	.datac(read_latency_shift_reg_0),
	.datad(\mem_used[0]~q ),
	.cin(gnd),
	.combout(\mem_used[1]~2_combout ),
	.cout());
defparam \mem_used[1]~2 .lut_mask = 16'hEFFF;
defparam \mem_used[1]~2 .sum_lutc_input = "datac";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclone10lp_lcell_comb \mem~0 (
	.dataa(\mem[1][74]~q ),
	.datab(saved_grant_1),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~0_combout ),
	.cout());
defparam \mem~0 .lut_mask = 16'hAACC;
defparam \mem~0 .sum_lutc_input = "datac";

dffeas \mem[1][56] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][56]~q ),
	.prn(vcc));
defparam \mem[1][56] .is_wysiwyg = "true";
defparam \mem[1][56] .power_up = "low";

cyclone10lp_lcell_comb \mem~1 (
	.dataa(\mem[1][56]~q ),
	.datab(src_data_56),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~1_combout ),
	.cout());
defparam \mem~1 .lut_mask = 16'hAACC;
defparam \mem~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \write~0 (
	.dataa(rst1),
	.datab(wait_latency_counter_1),
	.datac(src_valid),
	.datad(src_valid1),
	.cin(gnd),
	.combout(\write~0_combout ),
	.cout());
defparam \write~0 .lut_mask = 16'hFFFB;
defparam \write~0 .sum_lutc_input = "datac";

endmodule

module processor_altera_avalon_sc_fifo_6 (
	reset,
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	saved_grant_1,
	mem_used_1,
	cp_ready,
	cp_ready1,
	WideOr1,
	src_data_56,
	read_latency_shift_reg,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	read_latency_shift_reg_0;
output 	mem_74_0;
output 	mem_56_0;
input 	saved_grant_1;
output 	mem_used_1;
input 	cp_ready;
input 	cp_ready1;
input 	WideOr1;
input 	src_data_56;
input 	read_latency_shift_reg;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem[1][74]~q ;
wire \mem~0_combout ;
wire \mem_used[0]~3_combout ;
wire \mem_used[0]~4_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem[1][56]~q ;
wire \mem~1_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~2_combout ;


dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][56] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_56_0),
	.prn(vcc));
defparam \mem[0][56] .is_wysiwyg = "true";
defparam \mem[0][56] .power_up = "low";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclone10lp_lcell_comb \mem~0 (
	.dataa(\mem[1][74]~q ),
	.datab(saved_grant_1),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~0_combout ),
	.cout());
defparam \mem~0 .lut_mask = 16'hAACC;
defparam \mem~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_used[0]~3 (
	.dataa(\mem_used[0]~q ),
	.datab(mem_used_1),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hEEFF;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_used[0]~4 (
	.dataa(\mem_used[0]~3_combout ),
	.datab(WideOr1),
	.datac(src_data_56),
	.datad(cp_ready1),
	.cin(gnd),
	.combout(\mem_used[0]~4_combout ),
	.cout());
defparam \mem_used[0]~4 .lut_mask = 16'hFEFF;
defparam \mem_used[0]~4 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclone10lp_lcell_comb \mem_used[1]~0 (
	.dataa(\mem_used[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hFF55;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

dffeas \mem[1][56] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][56]~q ),
	.prn(vcc));
defparam \mem[1][56] .is_wysiwyg = "true";
defparam \mem[1][56] .power_up = "low";

cyclone10lp_lcell_comb \mem~1 (
	.dataa(\mem[1][56]~q ),
	.datab(src_data_56),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~1_combout ),
	.cout());
defparam \mem~1 .lut_mask = 16'hAACC;
defparam \mem~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_used[1]~1 (
	.dataa(mem_used_1),
	.datab(gnd),
	.datac(read_latency_shift_reg_0),
	.datad(\mem_used[0]~q ),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hAFFF;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_used[1]~2 (
	.dataa(\mem_used[1]~1_combout ),
	.datab(cp_ready),
	.datac(read_latency_shift_reg),
	.datad(\mem_used[1]~0_combout ),
	.cin(gnd),
	.combout(\mem_used[1]~2_combout ),
	.cout());
defparam \mem_used[1]~2 .lut_mask = 16'hFEFF;
defparam \mem_used[1]~2 .sum_lutc_input = "datac";

endmodule

module processor_altera_avalon_sc_fifo_7 (
	reset,
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	mem_used_1,
	uav_waitrequest,
	saved_grant_1,
	WideOr1,
	src_data_56,
	read_latency_shift_reg,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	read_latency_shift_reg_0;
output 	mem_74_0;
output 	mem_56_0;
output 	mem_used_1;
input 	uav_waitrequest;
input 	saved_grant_1;
input 	WideOr1;
input 	src_data_56;
input 	read_latency_shift_reg;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem[1][74]~q ;
wire \mem~0_combout ;
wire \mem_used[0]~3_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem[1][56]~q ;
wire \mem~1_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~2_combout ;


dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][56] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_56_0),
	.prn(vcc));
defparam \mem[0][56] .is_wysiwyg = "true";
defparam \mem[0][56] .power_up = "low";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclone10lp_lcell_comb \mem~0 (
	.dataa(\mem[1][74]~q ),
	.datab(saved_grant_1),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~0_combout ),
	.cout());
defparam \mem~0 .lut_mask = 16'hAACC;
defparam \mem~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_used[0]~3 (
	.dataa(read_latency_shift_reg),
	.datab(\mem_used[0]~q ),
	.datac(mem_used_1),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hFEFF;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclone10lp_lcell_comb \mem_used[1]~0 (
	.dataa(\mem_used[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hFF55;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

dffeas \mem[1][56] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][56]~q ),
	.prn(vcc));
defparam \mem[1][56] .is_wysiwyg = "true";
defparam \mem[1][56] .power_up = "low";

cyclone10lp_lcell_comb \mem~1 (
	.dataa(\mem[1][56]~q ),
	.datab(src_data_56),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~1_combout ),
	.cout());
defparam \mem~1 .lut_mask = 16'hAACC;
defparam \mem~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_used[1]~1 (
	.dataa(WideOr1),
	.datab(src_data_56),
	.datac(\mem_used[1]~0_combout ),
	.datad(uav_waitrequest),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hEFFF;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_used[1]~2 (
	.dataa(\mem_used[1]~1_combout ),
	.datab(mem_used_1),
	.datac(read_latency_shift_reg_0),
	.datad(\mem_used[0]~q ),
	.cin(gnd),
	.combout(\mem_used[1]~2_combout ),
	.cout());
defparam \mem_used[1]~2 .lut_mask = 16'hEFFF;
defparam \mem_used[1]~2 .sum_lutc_input = "datac";

endmodule

module processor_altera_merlin_master_agent (
	d_write,
	write_accepted,
	rst1,
	read_accepted,
	d_read,
	cp_valid,
	cp_valid1)/* synthesis synthesis_greybox=1 */;
input 	d_write;
input 	write_accepted;
input 	rst1;
input 	read_accepted;
input 	d_read;
output 	cp_valid;
output 	cp_valid1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclone10lp_lcell_comb \cp_valid~0 (
	.dataa(write_accepted),
	.datab(read_accepted),
	.datac(d_read),
	.datad(d_write),
	.cin(gnd),
	.combout(cp_valid),
	.cout());
defparam \cp_valid~0 .lut_mask = 16'hEFFF;
defparam \cp_valid~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \cp_valid~1 (
	.dataa(rst1),
	.datab(gnd),
	.datac(gnd),
	.datad(cp_valid),
	.cin(gnd),
	.combout(cp_valid1),
	.cout());
defparam \cp_valid~1 .lut_mask = 16'hAAFF;
defparam \cp_valid~1 .sum_lutc_input = "datac";

endmodule

module processor_altera_merlin_master_agent_1 (
	rst1,
	i_read,
	read_accepted,
	cp_valid1)/* synthesis synthesis_greybox=1 */;
input 	rst1;
input 	i_read;
input 	read_accepted;
output 	cp_valid1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclone10lp_lcell_comb cp_valid(
	.dataa(rst1),
	.datab(gnd),
	.datac(i_read),
	.datad(read_accepted),
	.cin(gnd),
	.combout(cp_valid1),
	.cout());
defparam cp_valid.lut_mask = 16'hAFFF;
defparam cp_valid.sum_lutc_input = "datac";

endmodule

module processor_altera_merlin_master_translator (
	reset,
	d_write,
	write_accepted1,
	rst1,
	read_accepted1,
	d_read,
	cp_valid,
	WideOr1,
	WideOr0,
	av_waitrequest,
	uav_read1,
	uav_write,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	d_write;
output 	write_accepted1;
input 	rst1;
output 	read_accepted1;
input 	d_read;
input 	cp_valid;
input 	WideOr1;
input 	WideOr0;
output 	av_waitrequest;
output 	uav_read1;
output 	uav_write;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_accepted~0_combout ;
wire \write_accepted~0_combout ;
wire \read_accepted~1_combout ;
wire \end_begintransfer~0_combout ;
wire \end_begintransfer~q ;
wire \av_waitrequest~0_combout ;


dffeas write_accepted(
	.clk(clk),
	.d(\write_accepted~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(write_accepted1),
	.prn(vcc));
defparam write_accepted.is_wysiwyg = "true";
defparam write_accepted.power_up = "low";

dffeas read_accepted(
	.clk(clk),
	.d(\read_accepted~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_accepted1),
	.prn(vcc));
defparam read_accepted.is_wysiwyg = "true";
defparam read_accepted.power_up = "low";

cyclone10lp_lcell_comb \av_waitrequest~1 (
	.dataa(d_read),
	.datab(WideOr1),
	.datac(d_write),
	.datad(\av_waitrequest~0_combout ),
	.cin(gnd),
	.combout(av_waitrequest),
	.cout());
defparam \av_waitrequest~1 .lut_mask = 16'h8DFF;
defparam \av_waitrequest~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb uav_read(
	.dataa(d_read),
	.datab(gnd),
	.datac(gnd),
	.datad(read_accepted1),
	.cin(gnd),
	.combout(uav_read1),
	.cout());
defparam uav_read.lut_mask = 16'hAAFF;
defparam uav_read.sum_lutc_input = "datac";

cyclone10lp_lcell_comb \uav_write~0 (
	.dataa(d_write),
	.datab(gnd),
	.datac(gnd),
	.datad(write_accepted1),
	.cin(gnd),
	.combout(uav_write),
	.cout());
defparam \uav_write~0 .lut_mask = 16'hAAFF;
defparam \uav_write~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \read_accepted~0 (
	.dataa(rst1),
	.datab(WideOr0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\read_accepted~0_combout ),
	.cout());
defparam \read_accepted~0 .lut_mask = 16'hEEEE;
defparam \read_accepted~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \write_accepted~0 (
	.dataa(av_waitrequest),
	.datab(write_accepted1),
	.datac(d_write),
	.datad(\read_accepted~0_combout ),
	.cin(gnd),
	.combout(\write_accepted~0_combout ),
	.cout());
defparam \write_accepted~0 .lut_mask = 16'hFFFE;
defparam \write_accepted~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \read_accepted~1 (
	.dataa(WideOr1),
	.datab(read_accepted1),
	.datac(d_read),
	.datad(\read_accepted~0_combout ),
	.cin(gnd),
	.combout(\read_accepted~1_combout ),
	.cout());
defparam \read_accepted~1 .lut_mask = 16'hFFFE;
defparam \read_accepted~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \end_begintransfer~0 (
	.dataa(\end_begintransfer~q ),
	.datab(cp_valid),
	.datac(rst1),
	.datad(WideOr0),
	.cin(gnd),
	.combout(\end_begintransfer~0_combout ),
	.cout());
defparam \end_begintransfer~0 .lut_mask = 16'hBFFF;
defparam \end_begintransfer~0 .sum_lutc_input = "datac";

dffeas end_begintransfer(
	.clk(clk),
	.d(\end_begintransfer~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\end_begintransfer~q ),
	.prn(vcc));
defparam end_begintransfer.is_wysiwyg = "true";
defparam end_begintransfer.power_up = "low";

cyclone10lp_lcell_comb \av_waitrequest~0 (
	.dataa(rst1),
	.datab(\end_begintransfer~q ),
	.datac(write_accepted1),
	.datad(WideOr0),
	.cin(gnd),
	.combout(\av_waitrequest~0_combout ),
	.cout());
defparam \av_waitrequest~0 .lut_mask = 16'hFFFE;
defparam \av_waitrequest~0 .sum_lutc_input = "datac";

endmodule

module processor_altera_merlin_master_translator_1 (
	reset,
	saved_grant_1,
	rst1,
	i_read,
	read_accepted1,
	Equal4,
	mem_used_1,
	saved_grant_11,
	mem_used_11,
	saved_grant_12,
	uav_read1,
	Equal6,
	cp_ready,
	mem_used_12,
	mem_used_13,
	uav_waitrequest,
	sink_ready,
	cp_ready1,
	saved_grant_13,
	WideOr1,
	WideOr11,
	Equal7,
	saved_grant_14,
	saved_grant_15,
	write,
	Equal1,
	saved_grant_16,
	Equal2,
	src_channel_2,
	saved_grant_17,
	Equal5,
	cp_ready2,
	Equal41,
	always1,
	cp_ready3,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	saved_grant_1;
input 	rst1;
input 	i_read;
output 	read_accepted1;
input 	Equal4;
input 	mem_used_1;
input 	saved_grant_11;
input 	mem_used_11;
input 	saved_grant_12;
output 	uav_read1;
input 	Equal6;
input 	cp_ready;
input 	mem_used_12;
input 	mem_used_13;
input 	uav_waitrequest;
input 	sink_ready;
input 	cp_ready1;
input 	saved_grant_13;
input 	WideOr1;
input 	WideOr11;
input 	Equal7;
input 	saved_grant_14;
input 	saved_grant_15;
input 	write;
input 	Equal1;
input 	saved_grant_16;
input 	Equal2;
input 	src_channel_2;
input 	saved_grant_17;
input 	Equal5;
input 	cp_ready2;
input 	Equal41;
input 	always1;
input 	cp_ready3;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_accepted~0_combout ;
wire \read_accepted~1_combout ;
wire \read_accepted~2_combout ;
wire \read_accepted~3_combout ;
wire \read_accepted~4_combout ;
wire \read_accepted~5_combout ;
wire \read_accepted~6_combout ;
wire \read_accepted~7_combout ;
wire \read_accepted~8_combout ;
wire \read_accepted~9_combout ;
wire \read_accepted~10_combout ;


dffeas read_accepted(
	.clk(clk),
	.d(\read_accepted~10_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_accepted1),
	.prn(vcc));
defparam read_accepted.is_wysiwyg = "true";
defparam read_accepted.power_up = "low";

cyclone10lp_lcell_comb uav_read(
	.dataa(gnd),
	.datab(gnd),
	.datac(i_read),
	.datad(read_accepted1),
	.cin(gnd),
	.combout(uav_read1),
	.cout());
defparam uav_read.lut_mask = 16'h0FFF;
defparam uav_read.sum_lutc_input = "datac";

cyclone10lp_lcell_comb \read_accepted~0 (
	.dataa(Equal4),
	.datab(Equal7),
	.datac(saved_grant_14),
	.datad(sink_ready),
	.cin(gnd),
	.combout(\read_accepted~0_combout ),
	.cout());
defparam \read_accepted~0 .lut_mask = 16'hFFFE;
defparam \read_accepted~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \read_accepted~1 (
	.dataa(\read_accepted~0_combout ),
	.datab(saved_grant_15),
	.datac(write),
	.datad(Equal1),
	.cin(gnd),
	.combout(\read_accepted~1_combout ),
	.cout());
defparam \read_accepted~1 .lut_mask = 16'hFEFF;
defparam \read_accepted~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \read_accepted~2 (
	.dataa(saved_grant_1),
	.datab(Equal6),
	.datac(cp_ready),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\read_accepted~2_combout ),
	.cout());
defparam \read_accepted~2 .lut_mask = 16'hFEFF;
defparam \read_accepted~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \read_accepted~3 (
	.dataa(saved_grant_16),
	.datab(mem_used_12),
	.datac(src_channel_2),
	.datad(gnd),
	.cin(gnd),
	.combout(\read_accepted~3_combout ),
	.cout());
defparam \read_accepted~3 .lut_mask = 16'hFBFB;
defparam \read_accepted~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \read_accepted~4 (
	.dataa(Equal2),
	.datab(saved_grant_17),
	.datac(mem_used_13),
	.datad(uav_waitrequest),
	.cin(gnd),
	.combout(\read_accepted~4_combout ),
	.cout());
defparam \read_accepted~4 .lut_mask = 16'hEFFF;
defparam \read_accepted~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \read_accepted~5 (
	.dataa(\read_accepted~4_combout ),
	.datab(saved_grant_12),
	.datac(Equal5),
	.datad(cp_ready2),
	.cin(gnd),
	.combout(\read_accepted~5_combout ),
	.cout());
defparam \read_accepted~5 .lut_mask = 16'hFEFF;
defparam \read_accepted~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \read_accepted~6 (
	.dataa(\read_accepted~1_combout ),
	.datab(\read_accepted~2_combout ),
	.datac(\read_accepted~3_combout ),
	.datad(\read_accepted~5_combout ),
	.cin(gnd),
	.combout(\read_accepted~6_combout ),
	.cout());
defparam \read_accepted~6 .lut_mask = 16'hFFFE;
defparam \read_accepted~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \read_accepted~7 (
	.dataa(saved_grant_11),
	.datab(Equal41),
	.datac(cp_ready1),
	.datad(mem_used_11),
	.cin(gnd),
	.combout(\read_accepted~7_combout ),
	.cout());
defparam \read_accepted~7 .lut_mask = 16'hFEFF;
defparam \read_accepted~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \read_accepted~8 (
	.dataa(\read_accepted~7_combout ),
	.datab(always1),
	.datac(saved_grant_13),
	.datad(cp_ready3),
	.cin(gnd),
	.combout(\read_accepted~8_combout ),
	.cout());
defparam \read_accepted~8 .lut_mask = 16'hFEFF;
defparam \read_accepted~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \read_accepted~9 (
	.dataa(rst1),
	.datab(i_read),
	.datac(\read_accepted~6_combout ),
	.datad(\read_accepted~8_combout ),
	.cin(gnd),
	.combout(\read_accepted~9_combout ),
	.cout());
defparam \read_accepted~9 .lut_mask = 16'hFFFB;
defparam \read_accepted~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \read_accepted~10 (
	.dataa(read_accepted1),
	.datab(WideOr1),
	.datac(WideOr11),
	.datad(\read_accepted~9_combout ),
	.cin(gnd),
	.combout(\read_accepted~10_combout ),
	.cout());
defparam \read_accepted~10 .lut_mask = 16'hFFBF;
defparam \read_accepted~10 .sum_lutc_input = "datac";

endmodule

module processor_altera_merlin_slave_agent_1 (
	rst1,
	always0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	cp_ready)/* synthesis synthesis_greybox=1 */;
input 	rst1;
input 	always0;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
output 	cp_ready;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclone10lp_lcell_comb \cp_ready~0 (
	.dataa(rst1),
	.datab(always0),
	.datac(wait_latency_counter_0),
	.datad(wait_latency_counter_1),
	.cin(gnd),
	.combout(cp_ready),
	.cout());
defparam \cp_ready~0 .lut_mask = 16'hBEFF;
defparam \cp_ready~0 .sum_lutc_input = "datac";

endmodule

module processor_altera_merlin_slave_agent_2 (
	WideOr1,
	mem,
	rf_source_valid)/* synthesis synthesis_greybox=1 */;
input 	WideOr1;
input 	mem;
output 	rf_source_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclone10lp_lcell_comb \rf_source_valid~0 (
	.dataa(WideOr1),
	.datab(mem),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(rf_source_valid),
	.cout());
defparam \rf_source_valid~0 .lut_mask = 16'hEEEE;
defparam \rf_source_valid~0 .sum_lutc_input = "datac";

endmodule

module processor_altera_merlin_slave_agent_4 (
	rst1,
	mem_used_1,
	always0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	cp_ready,
	cp_ready1)/* synthesis synthesis_greybox=1 */;
input 	rst1;
input 	mem_used_1;
input 	always0;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
output 	cp_ready;
output 	cp_ready1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \cp_ready~1_combout ;


cyclone10lp_lcell_comb \cp_ready~0 (
	.dataa(rst1),
	.datab(always0),
	.datac(wait_latency_counter_0),
	.datad(wait_latency_counter_1),
	.cin(gnd),
	.combout(cp_ready),
	.cout());
defparam \cp_ready~0 .lut_mask = 16'hBEFF;
defparam \cp_ready~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \cp_ready~2 (
	.dataa(mem_used_1),
	.datab(always0),
	.datac(wait_latency_counter_0),
	.datad(\cp_ready~1_combout ),
	.cin(gnd),
	.combout(cp_ready1),
	.cout());
defparam \cp_ready~2 .lut_mask = 16'hFFBE;
defparam \cp_ready~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \cp_ready~1 (
	.dataa(rst1),
	.datab(wait_latency_counter_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\cp_ready~1_combout ),
	.cout());
defparam \cp_ready~1 .lut_mask = 16'hDDDD;
defparam \cp_ready~1 .sum_lutc_input = "datac";

endmodule

module processor_altera_merlin_slave_agent_5 (
	rst1,
	always0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	cp_ready)/* synthesis synthesis_greybox=1 */;
input 	rst1;
input 	always0;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
output 	cp_ready;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclone10lp_lcell_comb \cp_ready~0 (
	.dataa(rst1),
	.datab(always0),
	.datac(wait_latency_counter_0),
	.datad(wait_latency_counter_1),
	.cin(gnd),
	.combout(cp_ready),
	.cout());
defparam \cp_ready~0 .lut_mask = 16'hBEFF;
defparam \cp_ready~0 .sum_lutc_input = "datac";

endmodule

module processor_altera_merlin_slave_agent_6 (
	d_write,
	write_accepted,
	rst1,
	saved_grant_0,
	wait_latency_counter_0,
	src_valid,
	src_valid1,
	mem_used_1,
	m0_write,
	wait_latency_counter_1,
	cp_ready1,
	cp_ready2)/* synthesis synthesis_greybox=1 */;
input 	d_write;
input 	write_accepted;
input 	rst1;
input 	saved_grant_0;
input 	wait_latency_counter_0;
input 	src_valid;
input 	src_valid1;
input 	mem_used_1;
output 	m0_write;
input 	wait_latency_counter_1;
output 	cp_ready1;
output 	cp_ready2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \m0_write~0_combout ;
wire \cp_ready~1_combout ;


cyclone10lp_lcell_comb \m0_write~1 (
	.dataa(\m0_write~0_combout ),
	.datab(src_valid),
	.datac(src_valid1),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(m0_write),
	.cout());
defparam \m0_write~1 .lut_mask = 16'hFEFF;
defparam \m0_write~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \cp_ready~0 (
	.dataa(rst1),
	.datab(wait_latency_counter_0),
	.datac(m0_write),
	.datad(wait_latency_counter_1),
	.cin(gnd),
	.combout(cp_ready1),
	.cout());
defparam \cp_ready~0 .lut_mask = 16'hBEFF;
defparam \cp_ready~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb cp_ready(
	.dataa(mem_used_1),
	.datab(wait_latency_counter_0),
	.datac(m0_write),
	.datad(\cp_ready~1_combout ),
	.cin(gnd),
	.combout(cp_ready2),
	.cout());
defparam cp_ready.lut_mask = 16'hFFBE;
defparam cp_ready.sum_lutc_input = "datac";

cyclone10lp_lcell_comb \m0_write~0 (
	.dataa(d_write),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\m0_write~0_combout ),
	.cout());
defparam \m0_write~0 .lut_mask = 16'hEEFF;
defparam \m0_write~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \cp_ready~1 (
	.dataa(rst1),
	.datab(wait_latency_counter_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\cp_ready~1_combout ),
	.cout());
defparam \cp_ready~1 .lut_mask = 16'hDDDD;
defparam \cp_ready~1 .sum_lutc_input = "datac";

endmodule

module processor_altera_merlin_slave_translator (
	av_readdata_pre_22,
	av_readdata_pre_16,
	av_readdata_pre_21,
	av_readdata_pre_20,
	av_readdata_pre_19,
	av_readdata_pre_18,
	av_readdata_pre_17,
	reset,
	rst1,
	read_latency_shift_reg_0,
	sink_ready,
	src_data_56,
	WideOr1,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_4,
	av_readdata_pre_3,
	av_readdata_pre_2,
	av_readdata_pre_5,
	av_readdata_pre_14,
	av_readdata_pre_15,
	av_readdata_pre_13,
	av_readdata_pre_12,
	av_readdata_pre_10,
	av_readdata_pre_9,
	av_readdata_pre_8,
	av_readdata_pre_7,
	av_readdata_pre_6,
	b_full,
	read_0,
	av_readdata,
	b_full1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_01,
	counter_reg_bit_51,
	counter_reg_bit_41,
	counter_reg_bit_31,
	counter_reg_bit_21,
	counter_reg_bit_11,
	clk)/* synthesis synthesis_greybox=1 */;
output 	av_readdata_pre_22;
output 	av_readdata_pre_16;
output 	av_readdata_pre_21;
output 	av_readdata_pre_20;
output 	av_readdata_pre_19;
output 	av_readdata_pre_18;
output 	av_readdata_pre_17;
input 	reset;
input 	rst1;
output 	read_latency_shift_reg_0;
input 	sink_ready;
input 	src_data_56;
input 	WideOr1;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_4;
output 	av_readdata_pre_3;
output 	av_readdata_pre_2;
output 	av_readdata_pre_5;
output 	av_readdata_pre_14;
output 	av_readdata_pre_15;
output 	av_readdata_pre_13;
output 	av_readdata_pre_12;
output 	av_readdata_pre_10;
output 	av_readdata_pre_9;
output 	av_readdata_pre_8;
output 	av_readdata_pre_7;
output 	av_readdata_pre_6;
input 	b_full;
input 	read_0;
input 	[31:0] av_readdata;
input 	b_full1;
input 	counter_reg_bit_5;
input 	counter_reg_bit_4;
input 	counter_reg_bit_3;
input 	counter_reg_bit_2;
input 	counter_reg_bit_1;
input 	counter_reg_bit_0;
input 	counter_reg_bit_01;
input 	counter_reg_bit_51;
input 	counter_reg_bit_41;
input 	counter_reg_bit_31;
input 	counter_reg_bit_21;
input 	counter_reg_bit_11;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \av_readdata_pre[16]~8 ;
wire \av_readdata_pre[17]~10 ;
wire \av_readdata_pre[18]~12 ;
wire \av_readdata_pre[19]~14 ;
wire \av_readdata_pre[20]~16 ;
wire \av_readdata_pre[21]~18 ;
wire \av_readdata_pre[22]~19_combout ;
wire \av_readdata_pre[16]~7_combout ;
wire \av_readdata_pre[21]~17_combout ;
wire \av_readdata_pre[20]~15_combout ;
wire \av_readdata_pre[19]~13_combout ;
wire \av_readdata_pre[18]~11_combout ;
wire \av_readdata_pre[17]~9_combout ;
wire \read_latency_shift_reg~0_combout ;
wire \av_readdata_pre[13]~21_combout ;


dffeas \av_readdata_pre[22] (
	.clk(clk),
	.d(\av_readdata_pre[22]~19_combout ),
	.asdata(b_full),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_22),
	.prn(vcc));
defparam \av_readdata_pre[22] .is_wysiwyg = "true";
defparam \av_readdata_pre[22] .power_up = "low";

dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(\av_readdata_pre[16]~7_combout ),
	.asdata(counter_reg_bit_01),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

dffeas \av_readdata_pre[21] (
	.clk(clk),
	.d(\av_readdata_pre[21]~17_combout ),
	.asdata(counter_reg_bit_51),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_21),
	.prn(vcc));
defparam \av_readdata_pre[21] .is_wysiwyg = "true";
defparam \av_readdata_pre[21] .power_up = "low";

dffeas \av_readdata_pre[20] (
	.clk(clk),
	.d(\av_readdata_pre[20]~15_combout ),
	.asdata(counter_reg_bit_41),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_20),
	.prn(vcc));
defparam \av_readdata_pre[20] .is_wysiwyg = "true";
defparam \av_readdata_pre[20] .power_up = "low";

dffeas \av_readdata_pre[19] (
	.clk(clk),
	.d(\av_readdata_pre[19]~13_combout ),
	.asdata(counter_reg_bit_31),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_19),
	.prn(vcc));
defparam \av_readdata_pre[19] .is_wysiwyg = "true";
defparam \av_readdata_pre[19] .power_up = "low";

dffeas \av_readdata_pre[18] (
	.clk(clk),
	.d(\av_readdata_pre[18]~11_combout ),
	.asdata(counter_reg_bit_21),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_18),
	.prn(vcc));
defparam \av_readdata_pre[18] .is_wysiwyg = "true";
defparam \av_readdata_pre[18] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(\av_readdata_pre[17]~9_combout ),
	.asdata(counter_reg_bit_11),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(\av_readdata_pre[13]~21_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

cyclone10lp_lcell_comb \av_readdata_pre[16]~7 (
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\av_readdata_pre[16]~7_combout ),
	.cout(\av_readdata_pre[16]~8 ));
defparam \av_readdata_pre[16]~7 .lut_mask = 16'hAA55;
defparam \av_readdata_pre[16]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_readdata_pre[17]~9 (
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\av_readdata_pre[16]~8 ),
	.combout(\av_readdata_pre[17]~9_combout ),
	.cout(\av_readdata_pre[17]~10 ));
defparam \av_readdata_pre[17]~9 .lut_mask = 16'h5AAF;
defparam \av_readdata_pre[17]~9 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \av_readdata_pre[18]~11 (
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\av_readdata_pre[17]~10 ),
	.combout(\av_readdata_pre[18]~11_combout ),
	.cout(\av_readdata_pre[18]~12 ));
defparam \av_readdata_pre[18]~11 .lut_mask = 16'h5A5F;
defparam \av_readdata_pre[18]~11 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \av_readdata_pre[19]~13 (
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\av_readdata_pre[18]~12 ),
	.combout(\av_readdata_pre[19]~13_combout ),
	.cout(\av_readdata_pre[19]~14 ));
defparam \av_readdata_pre[19]~13 .lut_mask = 16'h5AAF;
defparam \av_readdata_pre[19]~13 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \av_readdata_pre[20]~15 (
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\av_readdata_pre[19]~14 ),
	.combout(\av_readdata_pre[20]~15_combout ),
	.cout(\av_readdata_pre[20]~16 ));
defparam \av_readdata_pre[20]~15 .lut_mask = 16'h5A5F;
defparam \av_readdata_pre[20]~15 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \av_readdata_pre[21]~17 (
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\av_readdata_pre[20]~16 ),
	.combout(\av_readdata_pre[21]~17_combout ),
	.cout(\av_readdata_pre[21]~18 ));
defparam \av_readdata_pre[21]~17 .lut_mask = 16'h5AAF;
defparam \av_readdata_pre[21]~17 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \av_readdata_pre[22]~19 (
	.dataa(b_full1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\av_readdata_pre[21]~18 ),
	.combout(\av_readdata_pre[22]~19_combout ),
	.cout());
defparam \av_readdata_pre[22]~19 .lut_mask = 16'h5A5A;
defparam \av_readdata_pre[22]~19 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \read_latency_shift_reg~0 (
	.dataa(rst1),
	.datab(sink_ready),
	.datac(src_data_56),
	.datad(WideOr1),
	.cin(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hFFFE;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_readdata_pre[13]~21 (
	.dataa(b_full1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\av_readdata_pre[13]~21_combout ),
	.cout());
defparam \av_readdata_pre[13]~21 .lut_mask = 16'h5555;
defparam \av_readdata_pre[13]~21 .sum_lutc_input = "datac";

endmodule

module processor_altera_merlin_slave_translator_1 (
	reset,
	src_payload,
	rst1,
	mem_used_1,
	always0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	cp_ready,
	read_latency_shift_reg_0,
	WideOr1,
	src_data_56,
	read_latency_shift_reg,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	src_payload;
input 	rst1;
input 	mem_used_1;
input 	always0;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
input 	cp_ready;
output 	read_latency_shift_reg_0;
input 	WideOr1;
input 	src_data_56;
output 	read_latency_shift_reg;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter[0]~0_combout ;
wire \wait_latency_counter[0]~1_combout ;
wire \wait_latency_counter[0]~2_combout ;
wire \wait_latency_counter~3_combout ;
wire \wait_latency_counter~4_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(read_latency_shift_reg),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclone10lp_lcell_comb \read_latency_shift_reg~0 (
	.dataa(WideOr1),
	.datab(cp_ready),
	.datac(src_data_56),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(read_latency_shift_reg),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hFEFF;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

cyclone10lp_lcell_comb \wait_latency_counter[0]~0 (
	.dataa(rst1),
	.datab(src_payload),
	.datac(src_data_56),
	.datad(gnd),
	.cin(gnd),
	.combout(\wait_latency_counter[0]~0_combout ),
	.cout());
defparam \wait_latency_counter[0]~0 .lut_mask = 16'hFEFE;
defparam \wait_latency_counter[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wait_latency_counter[0]~1 (
	.dataa(gnd),
	.datab(always0),
	.datac(wait_latency_counter_0),
	.datad(wait_latency_counter_1),
	.cin(gnd),
	.combout(\wait_latency_counter[0]~1_combout ),
	.cout());
defparam \wait_latency_counter[0]~1 .lut_mask = 16'h3CFF;
defparam \wait_latency_counter[0]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wait_latency_counter[0]~2 (
	.dataa(WideOr1),
	.datab(\wait_latency_counter[0]~0_combout ),
	.datac(mem_used_1),
	.datad(\wait_latency_counter[0]~1_combout ),
	.cin(gnd),
	.combout(\wait_latency_counter[0]~2_combout ),
	.cout());
defparam \wait_latency_counter[0]~2 .lut_mask = 16'hEFFF;
defparam \wait_latency_counter[0]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wait_latency_counter~3 (
	.dataa(\wait_latency_counter[0]~2_combout ),
	.datab(gnd),
	.datac(wait_latency_counter_1),
	.datad(wait_latency_counter_0),
	.cin(gnd),
	.combout(\wait_latency_counter~3_combout ),
	.cout());
defparam \wait_latency_counter~3 .lut_mask = 16'hAFFA;
defparam \wait_latency_counter~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wait_latency_counter~4 (
	.dataa(wait_latency_counter_0),
	.datab(gnd),
	.datac(gnd),
	.datad(\wait_latency_counter[0]~2_combout ),
	.cin(gnd),
	.combout(\wait_latency_counter~4_combout ),
	.cout());
defparam \wait_latency_counter~4 .lut_mask = 16'hFF55;
defparam \wait_latency_counter~4 .sum_lutc_input = "datac";

endmodule

module processor_altera_merlin_slave_translator_2 (
	av_readdata,
	reset,
	rst1,
	read_latency_shift_reg_0,
	write,
	WideOr1,
	mem,
	av_readdata_pre_0,
	av_readdata_pre_22,
	av_readdata_pre_23,
	av_readdata_pre_24,
	av_readdata_pre_25,
	av_readdata_pre_26,
	av_readdata_pre_1,
	av_readdata_pre_4,
	av_readdata_pre_3,
	av_readdata_pre_2,
	av_readdata_pre_5,
	av_readdata_pre_14,
	av_readdata_pre_15,
	av_readdata_pre_11,
	av_readdata_pre_13,
	av_readdata_pre_16,
	av_readdata_pre_12,
	av_readdata_pre_10,
	av_readdata_pre_9,
	av_readdata_pre_8,
	av_readdata_pre_7,
	av_readdata_pre_6,
	av_readdata_pre_21,
	av_readdata_pre_20,
	av_readdata_pre_19,
	av_readdata_pre_18,
	av_readdata_pre_17,
	av_readdata_pre_27,
	av_readdata_pre_28,
	av_readdata_pre_29,
	av_readdata_pre_30,
	av_readdata_pre_31,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[31:0] av_readdata;
input 	reset;
input 	rst1;
output 	read_latency_shift_reg_0;
input 	write;
input 	WideOr1;
input 	mem;
output 	av_readdata_pre_0;
output 	av_readdata_pre_22;
output 	av_readdata_pre_23;
output 	av_readdata_pre_24;
output 	av_readdata_pre_25;
output 	av_readdata_pre_26;
output 	av_readdata_pre_1;
output 	av_readdata_pre_4;
output 	av_readdata_pre_3;
output 	av_readdata_pre_2;
output 	av_readdata_pre_5;
output 	av_readdata_pre_14;
output 	av_readdata_pre_15;
output 	av_readdata_pre_11;
output 	av_readdata_pre_13;
output 	av_readdata_pre_16;
output 	av_readdata_pre_12;
output 	av_readdata_pre_10;
output 	av_readdata_pre_9;
output 	av_readdata_pre_8;
output 	av_readdata_pre_7;
output 	av_readdata_pre_6;
output 	av_readdata_pre_21;
output 	av_readdata_pre_20;
output 	av_readdata_pre_19;
output 	av_readdata_pre_18;
output 	av_readdata_pre_17;
output 	av_readdata_pre_27;
output 	av_readdata_pre_28;
output 	av_readdata_pre_29;
output 	av_readdata_pre_30;
output 	av_readdata_pre_31;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[22] (
	.clk(clk),
	.d(av_readdata[22]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_22),
	.prn(vcc));
defparam \av_readdata_pre[22] .is_wysiwyg = "true";
defparam \av_readdata_pre[22] .power_up = "low";

dffeas \av_readdata_pre[23] (
	.clk(clk),
	.d(av_readdata[23]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_23),
	.prn(vcc));
defparam \av_readdata_pre[23] .is_wysiwyg = "true";
defparam \av_readdata_pre[23] .power_up = "low";

dffeas \av_readdata_pre[24] (
	.clk(clk),
	.d(av_readdata[24]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_24),
	.prn(vcc));
defparam \av_readdata_pre[24] .is_wysiwyg = "true";
defparam \av_readdata_pre[24] .power_up = "low";

dffeas \av_readdata_pre[25] (
	.clk(clk),
	.d(av_readdata[25]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_25),
	.prn(vcc));
defparam \av_readdata_pre[25] .is_wysiwyg = "true";
defparam \av_readdata_pre[25] .power_up = "low";

dffeas \av_readdata_pre[26] (
	.clk(clk),
	.d(av_readdata[26]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_26),
	.prn(vcc));
defparam \av_readdata_pre[26] .is_wysiwyg = "true";
defparam \av_readdata_pre[26] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[11] (
	.clk(clk),
	.d(av_readdata[11]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_11),
	.prn(vcc));
defparam \av_readdata_pre[11] .is_wysiwyg = "true";
defparam \av_readdata_pre[11] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(av_readdata[13]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(av_readdata[16]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[21] (
	.clk(clk),
	.d(av_readdata[21]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_21),
	.prn(vcc));
defparam \av_readdata_pre[21] .is_wysiwyg = "true";
defparam \av_readdata_pre[21] .power_up = "low";

dffeas \av_readdata_pre[20] (
	.clk(clk),
	.d(av_readdata[20]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_20),
	.prn(vcc));
defparam \av_readdata_pre[20] .is_wysiwyg = "true";
defparam \av_readdata_pre[20] .power_up = "low";

dffeas \av_readdata_pre[19] (
	.clk(clk),
	.d(av_readdata[19]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_19),
	.prn(vcc));
defparam \av_readdata_pre[19] .is_wysiwyg = "true";
defparam \av_readdata_pre[19] .power_up = "low";

dffeas \av_readdata_pre[18] (
	.clk(clk),
	.d(av_readdata[18]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_18),
	.prn(vcc));
defparam \av_readdata_pre[18] .is_wysiwyg = "true";
defparam \av_readdata_pre[18] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(av_readdata[17]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

dffeas \av_readdata_pre[27] (
	.clk(clk),
	.d(av_readdata[27]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_27),
	.prn(vcc));
defparam \av_readdata_pre[27] .is_wysiwyg = "true";
defparam \av_readdata_pre[27] .power_up = "low";

dffeas \av_readdata_pre[28] (
	.clk(clk),
	.d(av_readdata[28]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_28),
	.prn(vcc));
defparam \av_readdata_pre[28] .is_wysiwyg = "true";
defparam \av_readdata_pre[28] .power_up = "low";

dffeas \av_readdata_pre[29] (
	.clk(clk),
	.d(av_readdata[29]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_29),
	.prn(vcc));
defparam \av_readdata_pre[29] .is_wysiwyg = "true";
defparam \av_readdata_pre[29] .power_up = "low";

dffeas \av_readdata_pre[30] (
	.clk(clk),
	.d(av_readdata[30]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_30),
	.prn(vcc));
defparam \av_readdata_pre[30] .is_wysiwyg = "true";
defparam \av_readdata_pre[30] .power_up = "low";

dffeas \av_readdata_pre[31] (
	.clk(clk),
	.d(av_readdata[31]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_31),
	.prn(vcc));
defparam \av_readdata_pre[31] .is_wysiwyg = "true";
defparam \av_readdata_pre[31] .power_up = "low";

cyclone10lp_lcell_comb \read_latency_shift_reg~0 (
	.dataa(rst1),
	.datab(write),
	.datac(WideOr1),
	.datad(mem),
	.cin(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hFFFE;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

endmodule

module processor_altera_merlin_slave_translator_3 (
	reset,
	rst1,
	read_latency_shift_reg_0,
	mem_used_1,
	WideOr1,
	mem,
	read_latency_shift_reg,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	rst1;
output 	read_latency_shift_reg_0;
input 	mem_used_1;
input 	WideOr1;
input 	mem;
output 	read_latency_shift_reg;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(read_latency_shift_reg),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclone10lp_lcell_comb \read_latency_shift_reg~0 (
	.dataa(rst1),
	.datab(WideOr1),
	.datac(mem),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(read_latency_shift_reg),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hFEFF;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

endmodule

module processor_altera_merlin_slave_translator_4 (
	reset,
	rst1,
	saved_grant_0,
	src_valid,
	src_valid1,
	mem_used_1,
	always0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	cp_ready,
	uav_write,
	WideOr1,
	src_data_56,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	rst1;
input 	saved_grant_0;
input 	src_valid;
input 	src_valid1;
input 	mem_used_1;
input 	always0;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg_0;
input 	cp_ready;
input 	uav_write;
input 	WideOr1;
input 	src_data_56;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter[0]~0_combout ;
wire \wait_latency_counter[0]~1_combout ;
wire \wait_latency_counter~2_combout ;
wire \wait_latency_counter~3_combout ;
wire \read_latency_shift_reg~0_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

cyclone10lp_lcell_comb \wait_latency_counter[0]~0 (
	.dataa(rst1),
	.datab(src_data_56),
	.datac(uav_write),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(\wait_latency_counter[0]~0_combout ),
	.cout());
defparam \wait_latency_counter[0]~0 .lut_mask = 16'hFFFE;
defparam \wait_latency_counter[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wait_latency_counter[0]~1 (
	.dataa(\wait_latency_counter[0]~0_combout ),
	.datab(src_valid),
	.datac(src_valid1),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\wait_latency_counter[0]~1_combout ),
	.cout());
defparam \wait_latency_counter[0]~1 .lut_mask = 16'hFEFF;
defparam \wait_latency_counter[0]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wait_latency_counter~2 (
	.dataa(\wait_latency_counter[0]~1_combout ),
	.datab(always0),
	.datac(wait_latency_counter_1),
	.datad(wait_latency_counter_0),
	.cin(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.cout());
defparam \wait_latency_counter~2 .lut_mask = 16'hEFFE;
defparam \wait_latency_counter~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wait_latency_counter~3 (
	.dataa(wait_latency_counter_0),
	.datab(always0),
	.datac(wait_latency_counter_1),
	.datad(\wait_latency_counter[0]~1_combout ),
	.cin(gnd),
	.combout(\wait_latency_counter~3_combout ),
	.cout());
defparam \wait_latency_counter~3 .lut_mask = 16'hFFF7;
defparam \wait_latency_counter~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \read_latency_shift_reg~0 (
	.dataa(WideOr1),
	.datab(cp_ready),
	.datac(src_data_56),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hFEFF;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

endmodule

module processor_altera_merlin_slave_translator_5 (
	reset,
	rst1,
	saved_grant_0,
	src_valid,
	src_valid1,
	mem_used_1,
	always0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	cp_ready,
	WideOr1,
	src_data_56,
	uav_write,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_4,
	av_readdata_pre_3,
	av_readdata_pre_2,
	av_readdata_pre_5,
	av_readdata_pre_7,
	av_readdata_pre_6,
	av_readdata,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	rst1;
input 	saved_grant_0;
input 	src_valid;
input 	src_valid1;
input 	mem_used_1;
input 	always0;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg_0;
input 	cp_ready;
input 	WideOr1;
input 	src_data_56;
input 	uav_write;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_4;
output 	av_readdata_pre_3;
output 	av_readdata_pre_2;
output 	av_readdata_pre_5;
output 	av_readdata_pre_7;
output 	av_readdata_pre_6;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter[1]~0_combout ;
wire \wait_latency_counter[1]~1_combout ;
wire \wait_latency_counter~2_combout ;
wire \wait_latency_counter~3_combout ;
wire \read_latency_shift_reg~0_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

cyclone10lp_lcell_comb \wait_latency_counter[1]~0 (
	.dataa(rst1),
	.datab(src_data_56),
	.datac(uav_write),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(\wait_latency_counter[1]~0_combout ),
	.cout());
defparam \wait_latency_counter[1]~0 .lut_mask = 16'hFFFE;
defparam \wait_latency_counter[1]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wait_latency_counter[1]~1 (
	.dataa(\wait_latency_counter[1]~0_combout ),
	.datab(src_valid),
	.datac(src_valid1),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\wait_latency_counter[1]~1_combout ),
	.cout());
defparam \wait_latency_counter[1]~1 .lut_mask = 16'hFEFF;
defparam \wait_latency_counter[1]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wait_latency_counter~2 (
	.dataa(\wait_latency_counter[1]~1_combout ),
	.datab(always0),
	.datac(wait_latency_counter_1),
	.datad(wait_latency_counter_0),
	.cin(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.cout());
defparam \wait_latency_counter~2 .lut_mask = 16'hEFFE;
defparam \wait_latency_counter~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wait_latency_counter~3 (
	.dataa(wait_latency_counter_0),
	.datab(always0),
	.datac(wait_latency_counter_1),
	.datad(\wait_latency_counter[1]~1_combout ),
	.cin(gnd),
	.combout(\wait_latency_counter~3_combout ),
	.cout());
defparam \wait_latency_counter~3 .lut_mask = 16'hFFF7;
defparam \wait_latency_counter~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \read_latency_shift_reg~0 (
	.dataa(WideOr1),
	.datab(cp_ready),
	.datac(src_data_56),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hFEFF;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

endmodule

module processor_altera_merlin_slave_translator_6 (
	reset,
	rst1,
	read_latency_shift_reg_0,
	saved_grant_0,
	wait_latency_counter_0,
	src_valid,
	src_valid1,
	mem_used_1,
	m0_write,
	wait_latency_counter_1,
	cp_ready,
	uav_write,
	WideOr1,
	src_data_56,
	read_latency_shift_reg,
	av_readdata_pre_0,
	av_readdata,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	rst1;
output 	read_latency_shift_reg_0;
input 	saved_grant_0;
output 	wait_latency_counter_0;
input 	src_valid;
input 	src_valid1;
input 	mem_used_1;
input 	m0_write;
output 	wait_latency_counter_1;
input 	cp_ready;
input 	uav_write;
input 	WideOr1;
input 	src_data_56;
output 	read_latency_shift_reg;
output 	av_readdata_pre_0;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;
wire \wait_latency_counter[1]~0_combout ;
wire \wait_latency_counter[1]~1_combout ;
wire \wait_latency_counter~2_combout ;
wire \wait_latency_counter~3_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

cyclone10lp_lcell_comb \read_latency_shift_reg~1 (
	.dataa(src_data_56),
	.datab(src_valid),
	.datac(src_valid1),
	.datad(gnd),
	.cin(gnd),
	.combout(read_latency_shift_reg),
	.cout());
defparam \read_latency_shift_reg~1 .lut_mask = 16'hFEFE;
defparam \read_latency_shift_reg~1 .sum_lutc_input = "datac";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

cyclone10lp_lcell_comb \read_latency_shift_reg~0 (
	.dataa(WideOr1),
	.datab(cp_ready),
	.datac(src_data_56),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hFEFF;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wait_latency_counter[1]~0 (
	.dataa(rst1),
	.datab(src_data_56),
	.datac(uav_write),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(\wait_latency_counter[1]~0_combout ),
	.cout());
defparam \wait_latency_counter[1]~0 .lut_mask = 16'hFFFE;
defparam \wait_latency_counter[1]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wait_latency_counter[1]~1 (
	.dataa(\wait_latency_counter[1]~0_combout ),
	.datab(src_valid),
	.datac(src_valid1),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\wait_latency_counter[1]~1_combout ),
	.cout());
defparam \wait_latency_counter[1]~1 .lut_mask = 16'hFEFF;
defparam \wait_latency_counter[1]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wait_latency_counter~2 (
	.dataa(wait_latency_counter_0),
	.datab(m0_write),
	.datac(wait_latency_counter_1),
	.datad(\wait_latency_counter[1]~1_combout ),
	.cin(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.cout());
defparam \wait_latency_counter~2 .lut_mask = 16'hFFF7;
defparam \wait_latency_counter~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wait_latency_counter~3 (
	.dataa(\wait_latency_counter[1]~1_combout ),
	.datab(m0_write),
	.datac(wait_latency_counter_1),
	.datad(wait_latency_counter_0),
	.cin(gnd),
	.combout(\wait_latency_counter~3_combout ),
	.cout());
defparam \wait_latency_counter~3 .lut_mask = 16'hEFFE;
defparam \wait_latency_counter~3 .sum_lutc_input = "datac";

endmodule

module processor_altera_merlin_slave_translator_7 (
	reset,
	d_write,
	write_accepted,
	rst1,
	read_latency_shift_reg_0,
	saved_grant_0,
	mem_used_1,
	wait_latency_counter_1,
	uav_waitrequest,
	WideOr1,
	av_begintransfer,
	src_data_56,
	read_latency_shift_reg,
	rx_rd_strobe_onset,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_4,
	av_readdata_pre_3,
	av_readdata_pre_2,
	av_readdata_pre_5,
	av_readdata_pre_9,
	av_readdata_pre_8,
	av_readdata_pre_7,
	av_readdata_pre_6,
	av_readdata,
	end_begintransfer1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	d_write;
input 	write_accepted;
input 	rst1;
output 	read_latency_shift_reg_0;
input 	saved_grant_0;
input 	mem_used_1;
output 	wait_latency_counter_1;
output 	uav_waitrequest;
input 	WideOr1;
output 	av_begintransfer;
input 	src_data_56;
output 	read_latency_shift_reg;
input 	rx_rd_strobe_onset;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_4;
output 	av_readdata_pre_3;
output 	av_readdata_pre_2;
output 	av_readdata_pre_5;
output 	av_readdata_pre_9;
output 	av_readdata_pre_8;
output 	av_readdata_pre_7;
output 	av_readdata_pre_6;
input 	[31:0] av_readdata;
output 	end_begintransfer1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~2_combout ;
wire \wait_latency_counter~3_combout ;
wire \wait_latency_counter[0]~q ;
wire \wait_latency_counter~4_combout ;
wire \end_begintransfer~0_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(read_latency_shift_reg),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

cyclone10lp_lcell_comb \uav_waitrequest~0 (
	.dataa(wait_latency_counter_1),
	.datab(gnd),
	.datac(rst1),
	.datad(\wait_latency_counter[0]~q ),
	.cin(gnd),
	.combout(uav_waitrequest),
	.cout());
defparam \uav_waitrequest~0 .lut_mask = 16'hAFFF;
defparam \uav_waitrequest~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_begintransfer~0 (
	.dataa(d_write),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(write_accepted),
	.cin(gnd),
	.combout(av_begintransfer),
	.cout());
defparam \av_begintransfer~0 .lut_mask = 16'hEEFF;
defparam \av_begintransfer~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \read_latency_shift_reg~0 (
	.dataa(WideOr1),
	.datab(src_data_56),
	.datac(mem_used_1),
	.datad(uav_waitrequest),
	.cin(gnd),
	.combout(read_latency_shift_reg),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hEFFF;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas end_begintransfer(
	.clk(clk),
	.d(\end_begintransfer~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(end_begintransfer1),
	.prn(vcc));
defparam end_begintransfer.is_wysiwyg = "true";
defparam end_begintransfer.power_up = "low";

cyclone10lp_lcell_comb \wait_latency_counter~2 (
	.dataa(rst1),
	.datab(rx_rd_strobe_onset),
	.datac(av_begintransfer),
	.datad(src_data_56),
	.cin(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.cout());
defparam \wait_latency_counter~2 .lut_mask = 16'hFFFE;
defparam \wait_latency_counter~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wait_latency_counter~3 (
	.dataa(\wait_latency_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\wait_latency_counter~2_combout ),
	.cin(gnd),
	.combout(\wait_latency_counter~3_combout ),
	.cout());
defparam \wait_latency_counter~3 .lut_mask = 16'hFF55;
defparam \wait_latency_counter~3 .sum_lutc_input = "datac";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wait_latency_counter[0]~q ),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

cyclone10lp_lcell_comb \wait_latency_counter~4 (
	.dataa(wait_latency_counter_1),
	.datab(rst1),
	.datac(\wait_latency_counter[0]~q ),
	.datad(\wait_latency_counter~2_combout ),
	.cin(gnd),
	.combout(\wait_latency_counter~4_combout ),
	.cout());
defparam \wait_latency_counter~4 .lut_mask = 16'hFF7B;
defparam \wait_latency_counter~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \end_begintransfer~0 (
	.dataa(uav_waitrequest),
	.datab(\wait_latency_counter~2_combout ),
	.datac(end_begintransfer1),
	.datad(gnd),
	.cin(gnd),
	.combout(\end_begintransfer~0_combout ),
	.cout());
defparam \end_begintransfer~0 .lut_mask = 16'hFEFE;
defparam \end_begintransfer~0 .sum_lutc_input = "datac";

endmodule

module processor_processor_mm_interconnect_0_cmd_demux (
	W_alu_result_4,
	W_alu_result_5,
	W_alu_result_6,
	saved_grant_0,
	rst1,
	Equal4,
	mem_used_1,
	saved_grant_01,
	mem_used_11,
	saved_grant_02,
	mem_used_12,
	Equal6,
	cp_valid,
	cp_ready,
	Equal5,
	cp_ready1,
	Equal1,
	Equal7,
	Equal2,
	saved_grant_03,
	mem_used_13,
	always1,
	saved_grant_04,
	mem_used_14,
	uav_waitrequest,
	av_waitrequest,
	mem_used_15,
	sink_ready,
	saved_grant_05,
	saved_grant_06,
	waitrequest,
	mem_used_16,
	Equal41,
	cp_ready2,
	saved_grant_07,
	mem_used_17,
	cp_ready3,
	WideOr0,
	src2_valid)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	W_alu_result_5;
input 	W_alu_result_6;
input 	saved_grant_0;
input 	rst1;
input 	Equal4;
input 	mem_used_1;
input 	saved_grant_01;
input 	mem_used_11;
input 	saved_grant_02;
input 	mem_used_12;
input 	Equal6;
input 	cp_valid;
input 	cp_ready;
input 	Equal5;
input 	cp_ready1;
input 	Equal1;
input 	Equal7;
input 	Equal2;
input 	saved_grant_03;
input 	mem_used_13;
input 	always1;
input 	saved_grant_04;
input 	mem_used_14;
input 	uav_waitrequest;
input 	av_waitrequest;
input 	mem_used_15;
output 	sink_ready;
input 	saved_grant_05;
input 	saved_grant_06;
input 	waitrequest;
input 	mem_used_16;
input 	Equal41;
input 	cp_ready2;
input 	saved_grant_07;
input 	mem_used_17;
input 	cp_ready3;
output 	WideOr0;
output 	src2_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sink_ready~0_combout ;
wire \src2_valid~0_combout ;
wire \src2_valid~1_combout ;
wire \sink_ready~1_combout ;
wire \sink_ready~2_combout ;
wire \sink_ready~3_combout ;
wire \sink_ready~5_combout ;
wire \sink_ready~6_combout ;
wire \WideOr0~0_combout ;
wire \sink_ready~7_combout ;
wire \WideOr0~1_combout ;
wire \sink_ready~8_combout ;
wire \sink_ready~9_combout ;


cyclone10lp_lcell_comb \sink_ready~4 (
	.dataa(av_waitrequest),
	.datab(gnd),
	.datac(gnd),
	.datad(mem_used_15),
	.cin(gnd),
	.combout(sink_ready),
	.cout());
defparam \sink_ready~4 .lut_mask = 16'hAAFF;
defparam \sink_ready~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \WideOr0~2 (
	.dataa(\sink_ready~0_combout ),
	.datab(\WideOr0~1_combout ),
	.datac(\sink_ready~8_combout ),
	.datad(\sink_ready~9_combout ),
	.cin(gnd),
	.combout(WideOr0),
	.cout());
defparam \WideOr0~2 .lut_mask = 16'hFFFE;
defparam \WideOr0~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src2_valid~2 (
	.dataa(cp_valid),
	.datab(\src2_valid~0_combout ),
	.datac(\src2_valid~1_combout ),
	.datad(always1),
	.cin(gnd),
	.combout(src2_valid),
	.cout());
defparam \src2_valid~2 .lut_mask = 16'hFEFF;
defparam \src2_valid~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sink_ready~0 (
	.dataa(saved_grant_02),
	.datab(Equal5),
	.datac(cp_ready1),
	.datad(mem_used_12),
	.cin(gnd),
	.combout(\sink_ready~0_combout ),
	.cout());
defparam \sink_ready~0 .lut_mask = 16'hFEFF;
defparam \sink_ready~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src2_valid~0 (
	.dataa(W_alu_result_6),
	.datab(W_alu_result_4),
	.datac(W_alu_result_5),
	.datad(Equal4),
	.cin(gnd),
	.combout(\src2_valid~0_combout ),
	.cout());
defparam \src2_valid~0 .lut_mask = 16'hBFFF;
defparam \src2_valid~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src2_valid~1 (
	.dataa(Equal1),
	.datab(Equal4),
	.datac(Equal7),
	.datad(Equal2),
	.cin(gnd),
	.combout(\src2_valid~1_combout ),
	.cout());
defparam \src2_valid~1 .lut_mask = 16'hBFFF;
defparam \src2_valid~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sink_ready~1 (
	.dataa(rst1),
	.datab(saved_grant_03),
	.datac(gnd),
	.datad(mem_used_13),
	.cin(gnd),
	.combout(\sink_ready~1_combout ),
	.cout());
defparam \sink_ready~1 .lut_mask = 16'hEEFF;
defparam \sink_ready~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sink_ready~2 (
	.dataa(\src2_valid~0_combout ),
	.datab(\src2_valid~1_combout ),
	.datac(\sink_ready~1_combout ),
	.datad(always1),
	.cin(gnd),
	.combout(\sink_ready~2_combout ),
	.cout());
defparam \sink_ready~2 .lut_mask = 16'hFEFF;
defparam \sink_ready~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sink_ready~3 (
	.dataa(Equal2),
	.datab(saved_grant_04),
	.datac(mem_used_14),
	.datad(uav_waitrequest),
	.cin(gnd),
	.combout(\sink_ready~3_combout ),
	.cout());
defparam \sink_ready~3 .lut_mask = 16'hEFFF;
defparam \sink_ready~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sink_ready~5 (
	.dataa(Equal4),
	.datab(sink_ready),
	.datac(Equal7),
	.datad(saved_grant_05),
	.cin(gnd),
	.combout(\sink_ready~5_combout ),
	.cout());
defparam \sink_ready~5 .lut_mask = 16'hFFFE;
defparam \sink_ready~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sink_ready~6 (
	.dataa(saved_grant_06),
	.datab(waitrequest),
	.datac(mem_used_16),
	.datad(Equal1),
	.cin(gnd),
	.combout(\sink_ready~6_combout ),
	.cout());
defparam \sink_ready~6 .lut_mask = 16'hBFFF;
defparam \sink_ready~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \WideOr0~0 (
	.dataa(\sink_ready~2_combout ),
	.datab(\sink_ready~3_combout ),
	.datac(\sink_ready~5_combout ),
	.datad(\sink_ready~6_combout ),
	.cin(gnd),
	.combout(\WideOr0~0_combout ),
	.cout());
defparam \WideOr0~0 .lut_mask = 16'hFFFE;
defparam \WideOr0~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sink_ready~7 (
	.dataa(saved_grant_0),
	.datab(Equal6),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sink_ready~7_combout ),
	.cout());
defparam \sink_ready~7 .lut_mask = 16'hEEEE;
defparam \sink_ready~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \WideOr0~1 (
	.dataa(\WideOr0~0_combout ),
	.datab(cp_ready),
	.datac(\sink_ready~7_combout ),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\WideOr0~1_combout ),
	.cout());
defparam \WideOr0~1 .lut_mask = 16'hFEFF;
defparam \WideOr0~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sink_ready~8 (
	.dataa(saved_grant_01),
	.datab(Equal41),
	.datac(cp_ready2),
	.datad(mem_used_11),
	.cin(gnd),
	.combout(\sink_ready~8_combout ),
	.cout());
defparam \sink_ready~8 .lut_mask = 16'hFEFF;
defparam \sink_ready~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sink_ready~9 (
	.dataa(saved_grant_07),
	.datab(always1),
	.datac(cp_ready3),
	.datad(mem_used_17),
	.cin(gnd),
	.combout(\sink_ready~9_combout ),
	.cout());
defparam \sink_ready~9 .lut_mask = 16'hFEFF;
defparam \sink_ready~9 .sum_lutc_input = "datac";

endmodule

module processor_processor_mm_interconnect_0_cmd_demux_1 (
	rst1,
	i_read,
	read_accepted,
	cp_valid,
	Equal1,
	F_pc_10,
	F_pc_9,
	Equal4,
	F_pc_2,
	Equal41,
	uav_read,
	Equal6,
	Equal7,
	src_channel_2,
	Equal2,
	src_channel_21,
	Equal5,
	always1,
	src5_valid,
	src0_valid,
	src1_valid,
	src2_valid,
	src6_valid,
	src3_valid,
	src4_valid,
	src7_valid)/* synthesis synthesis_greybox=1 */;
input 	rst1;
input 	i_read;
input 	read_accepted;
input 	cp_valid;
input 	Equal1;
input 	F_pc_10;
input 	F_pc_9;
input 	Equal4;
input 	F_pc_2;
input 	Equal41;
input 	uav_read;
input 	Equal6;
input 	Equal7;
input 	src_channel_2;
input 	Equal2;
input 	src_channel_21;
input 	Equal5;
input 	always1;
output 	src5_valid;
output 	src0_valid;
output 	src1_valid;
output 	src2_valid;
output 	src6_valid;
output 	src3_valid;
output 	src4_valid;
output 	src7_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclone10lp_lcell_comb \src5_valid~0 (
	.dataa(rst1),
	.datab(uav_read),
	.datac(F_pc_2),
	.datad(Equal41),
	.cin(gnd),
	.combout(src5_valid),
	.cout());
defparam \src5_valid~0 .lut_mask = 16'hFFFE;
defparam \src5_valid~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src0_valid~0 (
	.dataa(rst1),
	.datab(uav_read),
	.datac(Equal4),
	.datad(Equal7),
	.cin(gnd),
	.combout(src0_valid),
	.cout());
defparam \src0_valid~0 .lut_mask = 16'hFFFE;
defparam \src0_valid~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src1_valid~0 (
	.dataa(cp_valid),
	.datab(Equal1),
	.datac(F_pc_9),
	.datad(F_pc_10),
	.cin(gnd),
	.combout(src1_valid),
	.cout());
defparam \src1_valid~0 .lut_mask = 16'hFEFF;
defparam \src1_valid~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src2_valid~0 (
	.dataa(cp_valid),
	.datab(src_channel_2),
	.datac(src_channel_21),
	.datad(always1),
	.cin(gnd),
	.combout(src2_valid),
	.cout());
defparam \src2_valid~0 .lut_mask = 16'hFEFF;
defparam \src2_valid~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src6_valid~0 (
	.dataa(rst1),
	.datab(uav_read),
	.datac(Equal41),
	.datad(F_pc_2),
	.cin(gnd),
	.combout(src6_valid),
	.cout());
defparam \src6_valid~0 .lut_mask = 16'hFEFF;
defparam \src6_valid~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src3_valid~2 (
	.dataa(i_read),
	.datab(read_accepted),
	.datac(rst1),
	.datad(Equal6),
	.cin(gnd),
	.combout(src3_valid),
	.cout());
defparam \src3_valid~2 .lut_mask = 16'hFFF7;
defparam \src3_valid~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src4_valid~2 (
	.dataa(i_read),
	.datab(read_accepted),
	.datac(rst1),
	.datad(Equal5),
	.cin(gnd),
	.combout(src4_valid),
	.cout());
defparam \src4_valid~2 .lut_mask = 16'hFFF7;
defparam \src4_valid~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src7_valid~2 (
	.dataa(i_read),
	.datab(read_accepted),
	.datac(rst1),
	.datad(Equal2),
	.cin(gnd),
	.combout(src7_valid),
	.cout());
defparam \src7_valid~2 .lut_mask = 16'hFFF7;
defparam \src7_valid~2 .sum_lutc_input = "datac";

endmodule

module processor_processor_mm_interconnect_0_cmd_mux (
	W_alu_result_2,
	d_writedata_0,
	r_sync_rst,
	rst1,
	Equal4,
	cp_valid,
	F_pc_0,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	uav_read,
	Equal7,
	sink_ready,
	saved_grant_0,
	saved_grant_1,
	uav_read1,
	src_data_56,
	src0_valid,
	WideOr11,
	src_data_38,
	src_payload,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_2;
input 	d_writedata_0;
input 	r_sync_rst;
input 	rst1;
input 	Equal4;
input 	cp_valid;
input 	F_pc_0;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
input 	uav_read;
input 	Equal7;
input 	sink_ready;
output 	saved_grant_0;
output 	saved_grant_1;
input 	uav_read1;
output 	src_data_56;
input 	src0_valid;
output 	WideOr11;
output 	src_data_38;
output 	src_payload;
output 	src_payload1;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
output 	src_payload7;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \update_grant~0_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~1_combout ;
wire \src_valid~2_combout ;


processor_altera_merlin_arbitrator_7 arb(
	.reset(r_sync_rst),
	.src0_valid(src0_valid),
	.grant_0(\arb|grant[0]~0_combout ),
	.update_grant(\update_grant~1_combout ),
	.grant_1(\arb|grant[1]~1_combout ),
	.src_valid(\src_valid~2_combout ),
	.clk(clk_clk));

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclone10lp_lcell_comb \src_data[56] (
	.dataa(uav_read),
	.datab(uav_read1),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_56),
	.cout());
defparam \src_data[56] .lut_mask = 16'hFFFE;
defparam \src_data[56] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb WideOr1(
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(\src_valid~2_combout ),
	.datad(src0_valid),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam WideOr1.lut_mask = 16'hFFFE;
defparam WideOr1.sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[38] (
	.dataa(W_alu_result_2),
	.datab(F_pc_0),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_38),
	.cout());
defparam \src_data[38] .lut_mask = 16'hFFFE;
defparam \src_data[38] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~0 (
	.dataa(d_writedata_7),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload),
	.cout());
defparam \src_payload~0 .lut_mask = 16'hEEEE;
defparam \src_payload~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~1 (
	.dataa(d_writedata_0),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload1),
	.cout());
defparam \src_payload~1 .lut_mask = 16'hEEEE;
defparam \src_payload~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~2 (
	.dataa(d_writedata_1),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload2),
	.cout());
defparam \src_payload~2 .lut_mask = 16'hEEEE;
defparam \src_payload~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~3 (
	.dataa(d_writedata_2),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload3),
	.cout());
defparam \src_payload~3 .lut_mask = 16'hEEEE;
defparam \src_payload~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~4 (
	.dataa(d_writedata_3),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload4),
	.cout());
defparam \src_payload~4 .lut_mask = 16'hEEEE;
defparam \src_payload~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~5 (
	.dataa(d_writedata_6),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload5),
	.cout());
defparam \src_payload~5 .lut_mask = 16'hEEEE;
defparam \src_payload~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~6 (
	.dataa(d_writedata_5),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload6),
	.cout());
defparam \src_payload~6 .lut_mask = 16'hEEEE;
defparam \src_payload~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~7 (
	.dataa(d_writedata_4),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload7),
	.cout());
defparam \src_payload~7 .lut_mask = 16'hEEEE;
defparam \src_payload~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \update_grant~0 (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\update_grant~0_combout ),
	.cout());
defparam \update_grant~0 .lut_mask = 16'hEEEE;
defparam \update_grant~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \packet_in_progress~0 (
	.dataa(\update_grant~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\packet_in_progress~0_combout ),
	.cout());
defparam \packet_in_progress~0 .lut_mask = 16'h5555;
defparam \packet_in_progress~0 .sum_lutc_input = "datac";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclone10lp_lcell_comb \update_grant~1 (
	.dataa(sink_ready),
	.datab(\update_grant~0_combout ),
	.datac(WideOr11),
	.datad(\packet_in_progress~q ),
	.cin(gnd),
	.combout(\update_grant~1_combout ),
	.cout());
defparam \update_grant~1 .lut_mask = 16'hACFF;
defparam \update_grant~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_valid~2 (
	.dataa(rst1),
	.datab(cp_valid),
	.datac(Equal4),
	.datad(Equal7),
	.cin(gnd),
	.combout(\src_valid~2_combout ),
	.cout());
defparam \src_valid~2 .lut_mask = 16'hFFFB;
defparam \src_valid~2 .sum_lutc_input = "datac";

endmodule

module processor_processor_mm_interconnect_0_cmd_mux_1 (
	W_alu_result_7,
	W_alu_result_10,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_4,
	W_alu_result_5,
	W_alu_result_6,
	W_alu_result_2,
	W_alu_result_3,
	d_writedata_24,
	d_writedata_25,
	d_writedata_26,
	d_writedata_27,
	d_writedata_28,
	d_writedata_29,
	d_writedata_30,
	d_writedata_31,
	d_writedata_0,
	r_sync_rst,
	rst1,
	F_pc_5,
	F_pc_8,
	F_pc_7,
	F_pc_6,
	F_pc_2,
	F_pc_3,
	F_pc_4,
	cp_valid,
	F_pc_1,
	F_pc_0,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	Equal1,
	saved_grant_0,
	waitrequest,
	mem_used_1,
	saved_grant_1,
	d_writedata_9,
	src1_valid,
	WideOr11,
	hbreak_enabled,
	src_data_46,
	d_byteenable_0,
	d_writedata_22,
	d_byteenable_2,
	d_writedata_23,
	d_byteenable_3,
	d_writedata_14,
	d_byteenable_1,
	d_writedata_15,
	d_writedata_11,
	d_writedata_13,
	d_writedata_16,
	d_writedata_12,
	d_writedata_10,
	d_writedata_8,
	d_writedata_21,
	d_writedata_20,
	d_writedata_19,
	d_writedata_18,
	d_writedata_17,
	src_payload,
	src_payload1,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_32,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_data_34,
	src_payload6,
	src_payload7,
	src_data_35,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_data_33,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_7;
input 	W_alu_result_10;
input 	W_alu_result_9;
input 	W_alu_result_8;
input 	W_alu_result_4;
input 	W_alu_result_5;
input 	W_alu_result_6;
input 	W_alu_result_2;
input 	W_alu_result_3;
input 	d_writedata_24;
input 	d_writedata_25;
input 	d_writedata_26;
input 	d_writedata_27;
input 	d_writedata_28;
input 	d_writedata_29;
input 	d_writedata_30;
input 	d_writedata_31;
input 	d_writedata_0;
input 	r_sync_rst;
input 	rst1;
input 	F_pc_5;
input 	F_pc_8;
input 	F_pc_7;
input 	F_pc_6;
input 	F_pc_2;
input 	F_pc_3;
input 	F_pc_4;
input 	cp_valid;
input 	F_pc_1;
input 	F_pc_0;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
input 	Equal1;
output 	saved_grant_0;
input 	waitrequest;
input 	mem_used_1;
output 	saved_grant_1;
input 	d_writedata_9;
input 	src1_valid;
output 	WideOr11;
input 	hbreak_enabled;
output 	src_data_46;
input 	d_byteenable_0;
input 	d_writedata_22;
input 	d_byteenable_2;
input 	d_writedata_23;
input 	d_byteenable_3;
input 	d_writedata_14;
input 	d_byteenable_1;
input 	d_writedata_15;
input 	d_writedata_11;
input 	d_writedata_13;
input 	d_writedata_16;
input 	d_writedata_12;
input 	d_writedata_10;
input 	d_writedata_8;
input 	d_writedata_21;
input 	d_writedata_20;
input 	d_writedata_19;
input 	d_writedata_18;
input 	d_writedata_17;
output 	src_payload;
output 	src_payload1;
output 	src_data_38;
output 	src_data_39;
output 	src_data_40;
output 	src_data_41;
output 	src_data_42;
output 	src_data_43;
output 	src_data_44;
output 	src_data_45;
output 	src_data_32;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_data_34;
output 	src_payload6;
output 	src_payload7;
output 	src_data_35;
output 	src_payload8;
output 	src_payload9;
output 	src_payload10;
output 	src_payload11;
output 	src_payload12;
output 	src_data_33;
output 	src_payload13;
output 	src_payload14;
output 	src_payload15;
output 	src_payload16;
output 	src_payload17;
output 	src_payload18;
output 	src_payload19;
output 	src_payload20;
output 	src_payload21;
output 	src_payload22;
output 	src_payload23;
output 	src_payload24;
output 	src_payload25;
output 	src_payload26;
output 	src_payload27;
output 	src_payload28;
output 	src_payload29;
output 	src_payload30;
output 	src_payload31;
output 	src_payload32;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \update_grant~0_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~1_combout ;
wire \src_valid~4_combout ;


processor_altera_merlin_arbitrator arb(
	.reset(r_sync_rst),
	.src1_valid(src1_valid),
	.grant_0(\arb|grant[0]~0_combout ),
	.update_grant(\update_grant~1_combout ),
	.grant_1(\arb|grant[1]~1_combout ),
	.src_valid(\src_valid~4_combout ),
	.clk(clk_clk));

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclone10lp_lcell_comb WideOr1(
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(\src_valid~4_combout ),
	.datad(src1_valid),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam WideOr1.lut_mask = 16'hFFFE;
defparam WideOr1.sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[46] (
	.dataa(F_pc_8),
	.datab(W_alu_result_10),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_46),
	.cout());
defparam \src_data[46] .lut_mask = 16'hFFFE;
defparam \src_data[46] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~0 (
	.dataa(saved_grant_0),
	.datab(hbreak_enabled),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload),
	.cout());
defparam \src_payload~0 .lut_mask = 16'hEEEE;
defparam \src_payload~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~1 (
	.dataa(d_writedata_0),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload1),
	.cout());
defparam \src_payload~1 .lut_mask = 16'hEEEE;
defparam \src_payload~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[38] (
	.dataa(W_alu_result_2),
	.datab(F_pc_0),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_38),
	.cout());
defparam \src_data[38] .lut_mask = 16'hFFFE;
defparam \src_data[38] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[39] (
	.dataa(W_alu_result_3),
	.datab(F_pc_1),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_39),
	.cout());
defparam \src_data[39] .lut_mask = 16'hFFFE;
defparam \src_data[39] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[40] (
	.dataa(F_pc_2),
	.datab(W_alu_result_4),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_40),
	.cout());
defparam \src_data[40] .lut_mask = 16'hFFFE;
defparam \src_data[40] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[41] (
	.dataa(F_pc_3),
	.datab(W_alu_result_5),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_41),
	.cout());
defparam \src_data[41] .lut_mask = 16'hFFFE;
defparam \src_data[41] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[42] (
	.dataa(F_pc_4),
	.datab(W_alu_result_6),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_42),
	.cout());
defparam \src_data[42] .lut_mask = 16'hFFFE;
defparam \src_data[42] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[43] (
	.dataa(F_pc_5),
	.datab(W_alu_result_7),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_43),
	.cout());
defparam \src_data[43] .lut_mask = 16'hFFFE;
defparam \src_data[43] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[44] (
	.dataa(F_pc_6),
	.datab(W_alu_result_8),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_44),
	.cout());
defparam \src_data[44] .lut_mask = 16'hFFFE;
defparam \src_data[44] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[45] (
	.dataa(F_pc_7),
	.datab(W_alu_result_9),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_45),
	.cout());
defparam \src_data[45] .lut_mask = 16'hFFFE;
defparam \src_data[45] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[32] (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(d_byteenable_0),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_32),
	.cout());
defparam \src_data[32] .lut_mask = 16'hFEFE;
defparam \src_data[32] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~2 (
	.dataa(d_writedata_1),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload2),
	.cout());
defparam \src_payload~2 .lut_mask = 16'hEEEE;
defparam \src_payload~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~3 (
	.dataa(d_writedata_3),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload3),
	.cout());
defparam \src_payload~3 .lut_mask = 16'hEEEE;
defparam \src_payload~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~4 (
	.dataa(d_writedata_2),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload4),
	.cout());
defparam \src_payload~4 .lut_mask = 16'hEEEE;
defparam \src_payload~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~5 (
	.dataa(saved_grant_0),
	.datab(d_writedata_22),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload5),
	.cout());
defparam \src_payload~5 .lut_mask = 16'hEEEE;
defparam \src_payload~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[34] (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(d_byteenable_2),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_34),
	.cout());
defparam \src_data[34] .lut_mask = 16'hFEFE;
defparam \src_data[34] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~6 (
	.dataa(saved_grant_0),
	.datab(d_writedata_23),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload6),
	.cout());
defparam \src_payload~6 .lut_mask = 16'hEEEE;
defparam \src_payload~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~7 (
	.dataa(saved_grant_0),
	.datab(d_writedata_24),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload7),
	.cout());
defparam \src_payload~7 .lut_mask = 16'hEEEE;
defparam \src_payload~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[35] (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(d_byteenable_3),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_35),
	.cout());
defparam \src_data[35] .lut_mask = 16'hFEFE;
defparam \src_data[35] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~8 (
	.dataa(saved_grant_0),
	.datab(d_writedata_25),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload8),
	.cout());
defparam \src_payload~8 .lut_mask = 16'hEEEE;
defparam \src_payload~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~9 (
	.dataa(saved_grant_0),
	.datab(d_writedata_26),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload9),
	.cout());
defparam \src_payload~9 .lut_mask = 16'hEEEE;
defparam \src_payload~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~10 (
	.dataa(d_writedata_4),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload10),
	.cout());
defparam \src_payload~10 .lut_mask = 16'hEEEE;
defparam \src_payload~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~11 (
	.dataa(d_writedata_5),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload11),
	.cout());
defparam \src_payload~11 .lut_mask = 16'hEEEE;
defparam \src_payload~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~12 (
	.dataa(saved_grant_0),
	.datab(d_writedata_14),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload12),
	.cout());
defparam \src_payload~12 .lut_mask = 16'hEEEE;
defparam \src_payload~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[33] (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(d_byteenable_1),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_33),
	.cout());
defparam \src_data[33] .lut_mask = 16'hFEFE;
defparam \src_data[33] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~13 (
	.dataa(saved_grant_0),
	.datab(d_writedata_15),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload13),
	.cout());
defparam \src_payload~13 .lut_mask = 16'hEEEE;
defparam \src_payload~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~14 (
	.dataa(saved_grant_0),
	.datab(d_writedata_11),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload14),
	.cout());
defparam \src_payload~14 .lut_mask = 16'hEEEE;
defparam \src_payload~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~15 (
	.dataa(saved_grant_0),
	.datab(d_writedata_13),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload15),
	.cout());
defparam \src_payload~15 .lut_mask = 16'hEEEE;
defparam \src_payload~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~16 (
	.dataa(saved_grant_0),
	.datab(d_writedata_16),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload16),
	.cout());
defparam \src_payload~16 .lut_mask = 16'hEEEE;
defparam \src_payload~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~17 (
	.dataa(saved_grant_0),
	.datab(d_writedata_12),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload17),
	.cout());
defparam \src_payload~17 .lut_mask = 16'hEEEE;
defparam \src_payload~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~18 (
	.dataa(saved_grant_0),
	.datab(d_writedata_10),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload18),
	.cout());
defparam \src_payload~18 .lut_mask = 16'hEEEE;
defparam \src_payload~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~19 (
	.dataa(saved_grant_0),
	.datab(d_writedata_9),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload19),
	.cout());
defparam \src_payload~19 .lut_mask = 16'hEEEE;
defparam \src_payload~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~20 (
	.dataa(saved_grant_0),
	.datab(d_writedata_8),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload20),
	.cout());
defparam \src_payload~20 .lut_mask = 16'hEEEE;
defparam \src_payload~20 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~21 (
	.dataa(d_writedata_7),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload21),
	.cout());
defparam \src_payload~21 .lut_mask = 16'hEEEE;
defparam \src_payload~21 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~22 (
	.dataa(d_writedata_6),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload22),
	.cout());
defparam \src_payload~22 .lut_mask = 16'hEEEE;
defparam \src_payload~22 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~23 (
	.dataa(saved_grant_0),
	.datab(d_writedata_21),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload23),
	.cout());
defparam \src_payload~23 .lut_mask = 16'hEEEE;
defparam \src_payload~23 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~24 (
	.dataa(saved_grant_0),
	.datab(d_writedata_20),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload24),
	.cout());
defparam \src_payload~24 .lut_mask = 16'hEEEE;
defparam \src_payload~24 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~25 (
	.dataa(saved_grant_0),
	.datab(d_writedata_19),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload25),
	.cout());
defparam \src_payload~25 .lut_mask = 16'hEEEE;
defparam \src_payload~25 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~26 (
	.dataa(saved_grant_0),
	.datab(d_writedata_18),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload26),
	.cout());
defparam \src_payload~26 .lut_mask = 16'hEEEE;
defparam \src_payload~26 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~27 (
	.dataa(saved_grant_0),
	.datab(d_writedata_17),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload27),
	.cout());
defparam \src_payload~27 .lut_mask = 16'hEEEE;
defparam \src_payload~27 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~28 (
	.dataa(saved_grant_0),
	.datab(d_writedata_27),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload28),
	.cout());
defparam \src_payload~28 .lut_mask = 16'hEEEE;
defparam \src_payload~28 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~29 (
	.dataa(saved_grant_0),
	.datab(d_writedata_28),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload29),
	.cout());
defparam \src_payload~29 .lut_mask = 16'hEEEE;
defparam \src_payload~29 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~30 (
	.dataa(saved_grant_0),
	.datab(d_writedata_29),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload30),
	.cout());
defparam \src_payload~30 .lut_mask = 16'hEEEE;
defparam \src_payload~30 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~31 (
	.dataa(saved_grant_0),
	.datab(d_writedata_30),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload31),
	.cout());
defparam \src_payload~31 .lut_mask = 16'hEEEE;
defparam \src_payload~31 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~32 (
	.dataa(saved_grant_0),
	.datab(d_writedata_31),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload32),
	.cout());
defparam \src_payload~32 .lut_mask = 16'hEEEE;
defparam \src_payload~32 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \update_grant~0 (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(waitrequest),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\update_grant~0_combout ),
	.cout());
defparam \update_grant~0 .lut_mask = 16'hEFFF;
defparam \update_grant~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \packet_in_progress~0 (
	.dataa(\update_grant~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\packet_in_progress~0_combout ),
	.cout());
defparam \packet_in_progress~0 .lut_mask = 16'h5555;
defparam \packet_in_progress~0 .sum_lutc_input = "datac";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclone10lp_lcell_comb \update_grant~1 (
	.dataa(\update_grant~0_combout ),
	.datab(WideOr11),
	.datac(gnd),
	.datad(\packet_in_progress~q ),
	.cin(gnd),
	.combout(\update_grant~1_combout ),
	.cout());
defparam \update_grant~1 .lut_mask = 16'h88BB;
defparam \update_grant~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_valid~4 (
	.dataa(rst1),
	.datab(cp_valid),
	.datac(Equal1),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_valid~4_combout ),
	.cout());
defparam \src_valid~4 .lut_mask = 16'hBFBF;
defparam \src_valid~4 .sum_lutc_input = "datac";

endmodule

module processor_altera_merlin_arbitrator (
	reset,
	src1_valid,
	grant_0,
	update_grant,
	grant_1,
	src_valid,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	src1_valid;
output 	grant_0;
input 	update_grant;
output 	grant_1;
input 	src_valid;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~q ;


cyclone10lp_lcell_comb \grant[0]~0 (
	.dataa(src_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(src1_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_0),
	.cout());
defparam \grant[0]~0 .lut_mask = 16'hEFFF;
defparam \grant[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \grant[1]~1 (
	.dataa(src1_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(src_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_1),
	.cout());
defparam \grant[1]~1 .lut_mask = 16'hEFFF;
defparam \grant[1]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \top_priority_reg[0]~0 (
	.dataa(update_grant),
	.datab(src1_valid),
	.datac(src_valid),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.cout());
defparam \top_priority_reg[0]~0 .lut_mask = 16'hFEFE;
defparam \top_priority_reg[0]~0 .sum_lutc_input = "datac";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cyclone10lp_lcell_comb \top_priority_reg[0]~1 (
	.dataa(grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.cout());
defparam \top_priority_reg[0]~1 .lut_mask = 16'h5555;
defparam \top_priority_reg[0]~1 .sum_lutc_input = "datac";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module processor_processor_mm_interconnect_0_cmd_mux_2 (
	W_alu_result_7,
	W_alu_result_14,
	W_alu_result_13,
	W_alu_result_12,
	W_alu_result_11,
	W_alu_result_10,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_4,
	W_alu_result_5,
	W_alu_result_6,
	W_alu_result_2,
	W_alu_result_3,
	d_writedata_24,
	d_writedata_25,
	d_writedata_26,
	d_writedata_27,
	d_writedata_28,
	d_writedata_29,
	d_writedata_30,
	d_writedata_31,
	d_writedata_0,
	r_sync_rst,
	rst1,
	F_pc_5,
	F_pc_12,
	F_pc_11,
	F_pc_10,
	F_pc_9,
	F_pc_8,
	F_pc_7,
	F_pc_6,
	F_pc_2,
	F_pc_3,
	F_pc_4,
	F_pc_1,
	F_pc_0,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	saved_grant_0,
	mem_used_1,
	saved_grant_1,
	d_writedata_9,
	src2_valid,
	src2_valid1,
	WideOr11,
	src_payload,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_46,
	src_data_47,
	src_data_48,
	src_data_49,
	src_data_50,
	d_byteenable_0,
	src_data_32,
	d_writedata_22,
	src_payload1,
	d_byteenable_2,
	src_data_34,
	d_writedata_23,
	src_payload2,
	src_payload3,
	d_byteenable_3,
	src_data_35,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	d_writedata_14,
	src_payload11,
	d_byteenable_1,
	src_data_33,
	d_writedata_15,
	src_payload12,
	d_writedata_11,
	src_payload13,
	d_writedata_13,
	src_payload14,
	d_writedata_16,
	src_payload15,
	d_writedata_12,
	src_payload16,
	d_writedata_10,
	src_payload17,
	src_payload18,
	d_writedata_8,
	src_payload19,
	src_payload20,
	src_payload21,
	d_writedata_21,
	src_payload22,
	d_writedata_20,
	src_payload23,
	d_writedata_19,
	src_payload24,
	d_writedata_18,
	src_payload25,
	d_writedata_17,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_7;
input 	W_alu_result_14;
input 	W_alu_result_13;
input 	W_alu_result_12;
input 	W_alu_result_11;
input 	W_alu_result_10;
input 	W_alu_result_9;
input 	W_alu_result_8;
input 	W_alu_result_4;
input 	W_alu_result_5;
input 	W_alu_result_6;
input 	W_alu_result_2;
input 	W_alu_result_3;
input 	d_writedata_24;
input 	d_writedata_25;
input 	d_writedata_26;
input 	d_writedata_27;
input 	d_writedata_28;
input 	d_writedata_29;
input 	d_writedata_30;
input 	d_writedata_31;
input 	d_writedata_0;
input 	r_sync_rst;
input 	rst1;
input 	F_pc_5;
input 	F_pc_12;
input 	F_pc_11;
input 	F_pc_10;
input 	F_pc_9;
input 	F_pc_8;
input 	F_pc_7;
input 	F_pc_6;
input 	F_pc_2;
input 	F_pc_3;
input 	F_pc_4;
input 	F_pc_1;
input 	F_pc_0;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
output 	saved_grant_0;
input 	mem_used_1;
output 	saved_grant_1;
input 	d_writedata_9;
input 	src2_valid;
input 	src2_valid1;
output 	WideOr11;
output 	src_payload;
output 	src_data_38;
output 	src_data_39;
output 	src_data_40;
output 	src_data_41;
output 	src_data_42;
output 	src_data_43;
output 	src_data_44;
output 	src_data_45;
output 	src_data_46;
output 	src_data_47;
output 	src_data_48;
output 	src_data_49;
output 	src_data_50;
input 	d_byteenable_0;
output 	src_data_32;
input 	d_writedata_22;
output 	src_payload1;
input 	d_byteenable_2;
output 	src_data_34;
input 	d_writedata_23;
output 	src_payload2;
output 	src_payload3;
input 	d_byteenable_3;
output 	src_data_35;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
output 	src_payload7;
output 	src_payload8;
output 	src_payload9;
output 	src_payload10;
input 	d_writedata_14;
output 	src_payload11;
input 	d_byteenable_1;
output 	src_data_33;
input 	d_writedata_15;
output 	src_payload12;
input 	d_writedata_11;
output 	src_payload13;
input 	d_writedata_13;
output 	src_payload14;
input 	d_writedata_16;
output 	src_payload15;
input 	d_writedata_12;
output 	src_payload16;
input 	d_writedata_10;
output 	src_payload17;
output 	src_payload18;
input 	d_writedata_8;
output 	src_payload19;
output 	src_payload20;
output 	src_payload21;
input 	d_writedata_21;
output 	src_payload22;
input 	d_writedata_20;
output 	src_payload23;
input 	d_writedata_19;
output 	src_payload24;
input 	d_writedata_18;
output 	src_payload25;
input 	d_writedata_17;
output 	src_payload26;
output 	src_payload27;
output 	src_payload28;
output 	src_payload29;
output 	src_payload30;
output 	src_payload31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \update_grant~0_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~1_combout ;


processor_altera_merlin_arbitrator_1 arb(
	.reset(r_sync_rst),
	.src2_valid(src2_valid),
	.src2_valid1(src2_valid1),
	.grant_0(\arb|grant[0]~0_combout ),
	.update_grant(\update_grant~1_combout ),
	.grant_1(\arb|grant[1]~1_combout ),
	.clk(clk_clk));

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclone10lp_lcell_comb WideOr1(
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(src2_valid),
	.datad(src2_valid1),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam WideOr1.lut_mask = 16'hFFFE;
defparam WideOr1.sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~0 (
	.dataa(d_writedata_0),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload),
	.cout());
defparam \src_payload~0 .lut_mask = 16'hEEEE;
defparam \src_payload~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[38] (
	.dataa(W_alu_result_2),
	.datab(F_pc_0),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_38),
	.cout());
defparam \src_data[38] .lut_mask = 16'hFFFE;
defparam \src_data[38] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[39] (
	.dataa(W_alu_result_3),
	.datab(F_pc_1),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_39),
	.cout());
defparam \src_data[39] .lut_mask = 16'hFFFE;
defparam \src_data[39] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[40] (
	.dataa(F_pc_2),
	.datab(W_alu_result_4),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_40),
	.cout());
defparam \src_data[40] .lut_mask = 16'hFFFE;
defparam \src_data[40] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[41] (
	.dataa(F_pc_3),
	.datab(W_alu_result_5),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_41),
	.cout());
defparam \src_data[41] .lut_mask = 16'hFFFE;
defparam \src_data[41] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[42] (
	.dataa(F_pc_4),
	.datab(W_alu_result_6),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_42),
	.cout());
defparam \src_data[42] .lut_mask = 16'hFFFE;
defparam \src_data[42] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[43] (
	.dataa(F_pc_5),
	.datab(W_alu_result_7),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_43),
	.cout());
defparam \src_data[43] .lut_mask = 16'hFFFE;
defparam \src_data[43] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[44] (
	.dataa(F_pc_6),
	.datab(W_alu_result_8),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_44),
	.cout());
defparam \src_data[44] .lut_mask = 16'hFFFE;
defparam \src_data[44] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[45] (
	.dataa(F_pc_7),
	.datab(W_alu_result_9),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_45),
	.cout());
defparam \src_data[45] .lut_mask = 16'hFFFE;
defparam \src_data[45] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[46] (
	.dataa(F_pc_8),
	.datab(W_alu_result_10),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_46),
	.cout());
defparam \src_data[46] .lut_mask = 16'hFFFE;
defparam \src_data[46] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[47] (
	.dataa(F_pc_9),
	.datab(W_alu_result_11),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_47),
	.cout());
defparam \src_data[47] .lut_mask = 16'hFFFE;
defparam \src_data[47] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[48] (
	.dataa(F_pc_10),
	.datab(W_alu_result_12),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_48),
	.cout());
defparam \src_data[48] .lut_mask = 16'hFFFE;
defparam \src_data[48] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[49] (
	.dataa(F_pc_11),
	.datab(W_alu_result_13),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_49),
	.cout());
defparam \src_data[49] .lut_mask = 16'hFFFE;
defparam \src_data[49] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[50] (
	.dataa(F_pc_12),
	.datab(W_alu_result_14),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_50),
	.cout());
defparam \src_data[50] .lut_mask = 16'hFFFE;
defparam \src_data[50] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[32] (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(d_byteenable_0),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_32),
	.cout());
defparam \src_data[32] .lut_mask = 16'hFEFE;
defparam \src_data[32] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~1 (
	.dataa(saved_grant_0),
	.datab(d_writedata_22),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload1),
	.cout());
defparam \src_payload~1 .lut_mask = 16'hEEEE;
defparam \src_payload~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[34] (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(d_byteenable_2),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_34),
	.cout());
defparam \src_data[34] .lut_mask = 16'hFEFE;
defparam \src_data[34] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~2 (
	.dataa(saved_grant_0),
	.datab(d_writedata_23),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload2),
	.cout());
defparam \src_payload~2 .lut_mask = 16'hEEEE;
defparam \src_payload~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~3 (
	.dataa(saved_grant_0),
	.datab(d_writedata_24),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload3),
	.cout());
defparam \src_payload~3 .lut_mask = 16'hEEEE;
defparam \src_payload~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[35] (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(d_byteenable_3),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_35),
	.cout());
defparam \src_data[35] .lut_mask = 16'hFEFE;
defparam \src_data[35] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~4 (
	.dataa(saved_grant_0),
	.datab(d_writedata_25),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload4),
	.cout());
defparam \src_payload~4 .lut_mask = 16'hEEEE;
defparam \src_payload~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~5 (
	.dataa(saved_grant_0),
	.datab(d_writedata_26),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload5),
	.cout());
defparam \src_payload~5 .lut_mask = 16'hEEEE;
defparam \src_payload~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~6 (
	.dataa(d_writedata_1),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload6),
	.cout());
defparam \src_payload~6 .lut_mask = 16'hEEEE;
defparam \src_payload~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~7 (
	.dataa(d_writedata_4),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload7),
	.cout());
defparam \src_payload~7 .lut_mask = 16'hEEEE;
defparam \src_payload~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~8 (
	.dataa(d_writedata_3),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload8),
	.cout());
defparam \src_payload~8 .lut_mask = 16'hEEEE;
defparam \src_payload~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~9 (
	.dataa(d_writedata_2),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload9),
	.cout());
defparam \src_payload~9 .lut_mask = 16'hEEEE;
defparam \src_payload~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~10 (
	.dataa(d_writedata_5),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload10),
	.cout());
defparam \src_payload~10 .lut_mask = 16'hEEEE;
defparam \src_payload~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~11 (
	.dataa(saved_grant_0),
	.datab(d_writedata_14),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload11),
	.cout());
defparam \src_payload~11 .lut_mask = 16'hEEEE;
defparam \src_payload~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[33] (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(d_byteenable_1),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_33),
	.cout());
defparam \src_data[33] .lut_mask = 16'hFEFE;
defparam \src_data[33] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~12 (
	.dataa(saved_grant_0),
	.datab(d_writedata_15),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload12),
	.cout());
defparam \src_payload~12 .lut_mask = 16'hEEEE;
defparam \src_payload~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~13 (
	.dataa(saved_grant_0),
	.datab(d_writedata_11),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload13),
	.cout());
defparam \src_payload~13 .lut_mask = 16'hEEEE;
defparam \src_payload~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~14 (
	.dataa(saved_grant_0),
	.datab(d_writedata_13),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload14),
	.cout());
defparam \src_payload~14 .lut_mask = 16'hEEEE;
defparam \src_payload~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~15 (
	.dataa(saved_grant_0),
	.datab(d_writedata_16),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload15),
	.cout());
defparam \src_payload~15 .lut_mask = 16'hEEEE;
defparam \src_payload~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~16 (
	.dataa(saved_grant_0),
	.datab(d_writedata_12),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload16),
	.cout());
defparam \src_payload~16 .lut_mask = 16'hEEEE;
defparam \src_payload~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~17 (
	.dataa(saved_grant_0),
	.datab(d_writedata_10),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload17),
	.cout());
defparam \src_payload~17 .lut_mask = 16'hEEEE;
defparam \src_payload~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~18 (
	.dataa(saved_grant_0),
	.datab(d_writedata_9),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload18),
	.cout());
defparam \src_payload~18 .lut_mask = 16'hEEEE;
defparam \src_payload~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~19 (
	.dataa(saved_grant_0),
	.datab(d_writedata_8),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload19),
	.cout());
defparam \src_payload~19 .lut_mask = 16'hEEEE;
defparam \src_payload~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~20 (
	.dataa(d_writedata_7),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload20),
	.cout());
defparam \src_payload~20 .lut_mask = 16'hEEEE;
defparam \src_payload~20 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~21 (
	.dataa(d_writedata_6),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload21),
	.cout());
defparam \src_payload~21 .lut_mask = 16'hEEEE;
defparam \src_payload~21 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~22 (
	.dataa(saved_grant_0),
	.datab(d_writedata_21),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload22),
	.cout());
defparam \src_payload~22 .lut_mask = 16'hEEEE;
defparam \src_payload~22 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~23 (
	.dataa(saved_grant_0),
	.datab(d_writedata_20),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload23),
	.cout());
defparam \src_payload~23 .lut_mask = 16'hEEEE;
defparam \src_payload~23 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~24 (
	.dataa(saved_grant_0),
	.datab(d_writedata_19),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload24),
	.cout());
defparam \src_payload~24 .lut_mask = 16'hEEEE;
defparam \src_payload~24 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~25 (
	.dataa(saved_grant_0),
	.datab(d_writedata_18),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload25),
	.cout());
defparam \src_payload~25 .lut_mask = 16'hEEEE;
defparam \src_payload~25 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~26 (
	.dataa(saved_grant_0),
	.datab(d_writedata_17),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload26),
	.cout());
defparam \src_payload~26 .lut_mask = 16'hEEEE;
defparam \src_payload~26 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~27 (
	.dataa(saved_grant_0),
	.datab(d_writedata_27),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload27),
	.cout());
defparam \src_payload~27 .lut_mask = 16'hEEEE;
defparam \src_payload~27 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~28 (
	.dataa(saved_grant_0),
	.datab(d_writedata_28),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload28),
	.cout());
defparam \src_payload~28 .lut_mask = 16'hEEEE;
defparam \src_payload~28 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~29 (
	.dataa(saved_grant_0),
	.datab(d_writedata_29),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload29),
	.cout());
defparam \src_payload~29 .lut_mask = 16'hEEEE;
defparam \src_payload~29 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~30 (
	.dataa(saved_grant_0),
	.datab(d_writedata_30),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload30),
	.cout());
defparam \src_payload~30 .lut_mask = 16'hEEEE;
defparam \src_payload~30 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~31 (
	.dataa(saved_grant_0),
	.datab(d_writedata_31),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload31),
	.cout());
defparam \src_payload~31 .lut_mask = 16'hEEEE;
defparam \src_payload~31 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \update_grant~0 (
	.dataa(rst1),
	.datab(saved_grant_1),
	.datac(saved_grant_0),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\update_grant~0_combout ),
	.cout());
defparam \update_grant~0 .lut_mask = 16'hFEFF;
defparam \update_grant~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \packet_in_progress~0 (
	.dataa(\update_grant~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\packet_in_progress~0_combout ),
	.cout());
defparam \packet_in_progress~0 .lut_mask = 16'h5555;
defparam \packet_in_progress~0 .sum_lutc_input = "datac";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclone10lp_lcell_comb \update_grant~1 (
	.dataa(\update_grant~0_combout ),
	.datab(WideOr11),
	.datac(gnd),
	.datad(\packet_in_progress~q ),
	.cin(gnd),
	.combout(\update_grant~1_combout ),
	.cout());
defparam \update_grant~1 .lut_mask = 16'h88BB;
defparam \update_grant~1 .sum_lutc_input = "datac";

endmodule

module processor_altera_merlin_arbitrator_1 (
	reset,
	src2_valid,
	src2_valid1,
	grant_0,
	update_grant,
	grant_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	src2_valid;
input 	src2_valid1;
output 	grant_0;
input 	update_grant;
output 	grant_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~q ;


cyclone10lp_lcell_comb \grant[0]~0 (
	.dataa(src2_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(src2_valid1),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_0),
	.cout());
defparam \grant[0]~0 .lut_mask = 16'hEFFF;
defparam \grant[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \grant[1]~1 (
	.dataa(src2_valid1),
	.datab(\top_priority_reg[1]~q ),
	.datac(src2_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_1),
	.cout());
defparam \grant[1]~1 .lut_mask = 16'hEFFF;
defparam \grant[1]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \top_priority_reg[0]~0 (
	.dataa(update_grant),
	.datab(src2_valid),
	.datac(src2_valid1),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.cout());
defparam \top_priority_reg[0]~0 .lut_mask = 16'hFEFE;
defparam \top_priority_reg[0]~0 .sum_lutc_input = "datac";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cyclone10lp_lcell_comb \top_priority_reg[0]~1 (
	.dataa(grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.cout());
defparam \top_priority_reg[0]~1 .lut_mask = 16'h5555;
defparam \top_priority_reg[0]~1 .sum_lutc_input = "datac";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module processor_processor_mm_interconnect_0_cmd_mux_3 (
	W_alu_result_4,
	W_alu_result_5,
	W_alu_result_6,
	r_sync_rst,
	saved_grant_0,
	d_write,
	write_accepted,
	src_payload,
	saved_grant_1,
	rst1,
	cp_valid,
	Equal4,
	F_pc_2,
	F_pc_3,
	F_pc_4,
	src_valid,
	Equal41,
	cp_valid1,
	src_valid1,
	mem_used_1,
	Equal6,
	uav_read,
	cp_ready,
	WideOr11,
	uav_read1,
	src_data_56,
	src3_valid,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	W_alu_result_5;
input 	W_alu_result_6;
input 	r_sync_rst;
output 	saved_grant_0;
input 	d_write;
input 	write_accepted;
output 	src_payload;
output 	saved_grant_1;
input 	rst1;
input 	cp_valid;
input 	Equal4;
input 	F_pc_2;
input 	F_pc_3;
input 	F_pc_4;
output 	src_valid;
input 	Equal41;
input 	cp_valid1;
output 	src_valid1;
input 	mem_used_1;
input 	Equal6;
input 	uav_read;
input 	cp_ready;
output 	WideOr11;
input 	uav_read1;
output 	src_data_56;
input 	src3_valid;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \src_valid~6_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;
wire \update_grant~1_combout ;
wire \src_valid~2_combout ;
wire \src_valid~4_combout ;


processor_altera_merlin_arbitrator_2 arb(
	.reset(r_sync_rst),
	.grant_0(\arb|grant[0]~0_combout ),
	.update_grant(\update_grant~1_combout ),
	.grant_1(\arb|grant[1]~1_combout ),
	.src_valid(\src_valid~6_combout ),
	.src3_valid(src3_valid),
	.clk(clk_clk));

cyclone10lp_lcell_comb \src_valid~6 (
	.dataa(rst1),
	.datab(cp_valid1),
	.datac(Equal6),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_valid~6_combout ),
	.cout());
defparam \src_valid~6 .lut_mask = 16'hFBFB;
defparam \src_valid~6 .sum_lutc_input = "datac";

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

cyclone10lp_lcell_comb \src_payload~0 (
	.dataa(saved_grant_0),
	.datab(d_write),
	.datac(gnd),
	.datad(write_accepted),
	.cin(gnd),
	.combout(src_payload),
	.cout());
defparam \src_payload~0 .lut_mask = 16'hEEFF;
defparam \src_payload~0 .sum_lutc_input = "datac";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclone10lp_lcell_comb \src_valid~3 (
	.dataa(saved_grant_1),
	.datab(cp_valid),
	.datac(Equal4),
	.datad(\src_valid~2_combout ),
	.cin(gnd),
	.combout(src_valid),
	.cout());
defparam \src_valid~3 .lut_mask = 16'hFFFE;
defparam \src_valid~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_valid~5 (
	.dataa(Equal41),
	.datab(rst1),
	.datac(cp_valid1),
	.datad(\src_valid~4_combout ),
	.cin(gnd),
	.combout(src_valid1),
	.cout());
defparam \src_valid~5 .lut_mask = 16'hFFEF;
defparam \src_valid~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb WideOr1(
	.dataa(src_valid),
	.datab(src_valid1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam WideOr1.lut_mask = 16'hEEEE;
defparam WideOr1.sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[56] (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(uav_read1),
	.datad(uav_read),
	.cin(gnd),
	.combout(src_data_56),
	.cout());
defparam \src_data[56] .lut_mask = 16'hFFFE;
defparam \src_data[56] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \packet_in_progress~0 (
	.dataa(\update_grant~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\packet_in_progress~0_combout ),
	.cout());
defparam \packet_in_progress~0 .lut_mask = 16'h5555;
defparam \packet_in_progress~0 .sum_lutc_input = "datac";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclone10lp_lcell_comb \update_grant~0 (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(cp_ready),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\update_grant~0_combout ),
	.cout());
defparam \update_grant~0 .lut_mask = 16'hFEFF;
defparam \update_grant~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \update_grant~1 (
	.dataa(src_valid),
	.datab(src_valid1),
	.datac(\packet_in_progress~q ),
	.datad(\update_grant~0_combout ),
	.cin(gnd),
	.combout(\update_grant~1_combout ),
	.cout());
defparam \update_grant~1 .lut_mask = 16'hFF6F;
defparam \update_grant~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_valid~2 (
	.dataa(F_pc_2),
	.datab(F_pc_3),
	.datac(F_pc_4),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_valid~2_combout ),
	.cout());
defparam \src_valid~2 .lut_mask = 16'hEFEF;
defparam \src_valid~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_valid~4 (
	.dataa(saved_grant_0),
	.datab(W_alu_result_4),
	.datac(W_alu_result_5),
	.datad(W_alu_result_6),
	.cin(gnd),
	.combout(\src_valid~4_combout ),
	.cout());
defparam \src_valid~4 .lut_mask = 16'hFEFF;
defparam \src_valid~4 .sum_lutc_input = "datac";

endmodule

module processor_altera_merlin_arbitrator_2 (
	reset,
	grant_0,
	update_grant,
	grant_1,
	src_valid,
	src3_valid,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
output 	grant_0;
input 	update_grant;
output 	grant_1;
input 	src_valid;
input 	src3_valid;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~q ;


cyclone10lp_lcell_comb \grant[0]~0 (
	.dataa(src_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(src3_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_0),
	.cout());
defparam \grant[0]~0 .lut_mask = 16'hEFFF;
defparam \grant[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \grant[1]~1 (
	.dataa(src3_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(src_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_1),
	.cout());
defparam \grant[1]~1 .lut_mask = 16'hEFFF;
defparam \grant[1]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \top_priority_reg[0]~0 (
	.dataa(update_grant),
	.datab(src3_valid),
	.datac(src_valid),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.cout());
defparam \top_priority_reg[0]~0 .lut_mask = 16'hFEFE;
defparam \top_priority_reg[0]~0 .sum_lutc_input = "datac";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cyclone10lp_lcell_comb \top_priority_reg[0]~1 (
	.dataa(grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.cout());
defparam \top_priority_reg[0]~1 .lut_mask = 16'h5555;
defparam \top_priority_reg[0]~1 .sum_lutc_input = "datac";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module processor_processor_mm_interconnect_0_cmd_mux_4 (
	W_alu_result_4,
	W_alu_result_5,
	W_alu_result_6,
	r_sync_rst,
	d_write,
	write_accepted,
	rst1,
	cp_valid,
	Equal4,
	F_pc_2,
	F_pc_3,
	F_pc_4,
	Equal41,
	cp_valid1,
	saved_grant_0,
	src_payload,
	saved_grant_1,
	src_valid,
	src_valid1,
	uav_read,
	Equal5,
	cp_ready,
	uav_read1,
	WideOr11,
	src_data_56,
	src_valid2,
	src4_valid,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	W_alu_result_5;
input 	W_alu_result_6;
input 	r_sync_rst;
input 	d_write;
input 	write_accepted;
input 	rst1;
input 	cp_valid;
input 	Equal4;
input 	F_pc_2;
input 	F_pc_3;
input 	F_pc_4;
input 	Equal41;
input 	cp_valid1;
output 	saved_grant_0;
output 	src_payload;
output 	saved_grant_1;
output 	src_valid;
output 	src_valid1;
input 	uav_read;
input 	Equal5;
input 	cp_ready;
input 	uav_read1;
output 	WideOr11;
output 	src_data_56;
output 	src_valid2;
input 	src4_valid;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \update_grant~0_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~1_combout ;
wire \src_valid~2_combout ;
wire \src_valid~4_combout ;


processor_altera_merlin_arbitrator_3 arb(
	.reset(r_sync_rst),
	.grant_0(\arb|grant[0]~0_combout ),
	.update_grant(\update_grant~1_combout ),
	.grant_1(\arb|grant[1]~1_combout ),
	.src_valid(src_valid2),
	.src4_valid(src4_valid),
	.clk(clk_clk));

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

cyclone10lp_lcell_comb \src_payload~0 (
	.dataa(d_write),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(write_accepted),
	.cin(gnd),
	.combout(src_payload),
	.cout());
defparam \src_payload~0 .lut_mask = 16'hEEFF;
defparam \src_payload~0 .sum_lutc_input = "datac";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclone10lp_lcell_comb \src_valid~3 (
	.dataa(cp_valid),
	.datab(F_pc_3),
	.datac(Equal4),
	.datad(\src_valid~2_combout ),
	.cin(gnd),
	.combout(src_valid),
	.cout());
defparam \src_valid~3 .lut_mask = 16'hFFFE;
defparam \src_valid~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_valid~5 (
	.dataa(saved_grant_0),
	.datab(cp_valid1),
	.datac(Equal41),
	.datad(\src_valid~4_combout ),
	.cin(gnd),
	.combout(src_valid1),
	.cout());
defparam \src_valid~5 .lut_mask = 16'hFFFB;
defparam \src_valid~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb WideOr1(
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(src_valid2),
	.datad(src4_valid),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam WideOr1.lut_mask = 16'hFFFE;
defparam WideOr1.sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[56] (
	.dataa(uav_read),
	.datab(uav_read1),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_56),
	.cout());
defparam \src_data[56] .lut_mask = 16'hFFFE;
defparam \src_data[56] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_valid~6 (
	.dataa(rst1),
	.datab(cp_valid1),
	.datac(Equal5),
	.datad(gnd),
	.cin(gnd),
	.combout(src_valid2),
	.cout());
defparam \src_valid~6 .lut_mask = 16'hFBFB;
defparam \src_valid~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \update_grant~0 (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\update_grant~0_combout ),
	.cout());
defparam \update_grant~0 .lut_mask = 16'hEEEE;
defparam \update_grant~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \packet_in_progress~0 (
	.dataa(\update_grant~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\packet_in_progress~0_combout ),
	.cout());
defparam \packet_in_progress~0 .lut_mask = 16'h5555;
defparam \packet_in_progress~0 .sum_lutc_input = "datac";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclone10lp_lcell_comb \update_grant~1 (
	.dataa(\update_grant~0_combout ),
	.datab(WideOr11),
	.datac(\packet_in_progress~q ),
	.datad(cp_ready),
	.cin(gnd),
	.combout(\update_grant~1_combout ),
	.cout());
defparam \update_grant~1 .lut_mask = 16'h8BFF;
defparam \update_grant~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_valid~2 (
	.dataa(saved_grant_1),
	.datab(F_pc_2),
	.datac(F_pc_4),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_valid~2_combout ),
	.cout());
defparam \src_valid~2 .lut_mask = 16'hBFBF;
defparam \src_valid~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_valid~4 (
	.dataa(rst1),
	.datab(W_alu_result_5),
	.datac(W_alu_result_4),
	.datad(W_alu_result_6),
	.cin(gnd),
	.combout(\src_valid~4_combout ),
	.cout());
defparam \src_valid~4 .lut_mask = 16'hEFFF;
defparam \src_valid~4 .sum_lutc_input = "datac";

endmodule

module processor_altera_merlin_arbitrator_3 (
	reset,
	grant_0,
	update_grant,
	grant_1,
	src_valid,
	src4_valid,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
output 	grant_0;
input 	update_grant;
output 	grant_1;
input 	src_valid;
input 	src4_valid;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~q ;


cyclone10lp_lcell_comb \grant[0]~0 (
	.dataa(src_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(src4_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_0),
	.cout());
defparam \grant[0]~0 .lut_mask = 16'hEFFF;
defparam \grant[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \grant[1]~1 (
	.dataa(src4_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(src_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_1),
	.cout());
defparam \grant[1]~1 .lut_mask = 16'hEFFF;
defparam \grant[1]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \top_priority_reg[0]~0 (
	.dataa(update_grant),
	.datab(src4_valid),
	.datac(src_valid),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.cout());
defparam \top_priority_reg[0]~0 .lut_mask = 16'hFEFE;
defparam \top_priority_reg[0]~0 .sum_lutc_input = "datac";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cyclone10lp_lcell_comb \top_priority_reg[0]~1 (
	.dataa(grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.cout());
defparam \top_priority_reg[0]~1 .lut_mask = 16'h5555;
defparam \top_priority_reg[0]~1 .sum_lutc_input = "datac";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module processor_processor_mm_interconnect_0_cmd_mux_5 (
	W_alu_result_4,
	W_alu_result_5,
	W_alu_result_6,
	r_sync_rst,
	d_write,
	write_accepted,
	rst1,
	cp_valid,
	F_pc_2,
	Equal4,
	cp_valid1,
	saved_grant_0,
	src_payload,
	saved_grant_1,
	Equal41,
	src_valid,
	src_valid1,
	uav_read,
	Equal42,
	uav_read1,
	src5_valid,
	write,
	WideOr11,
	src_data_56,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	W_alu_result_5;
input 	W_alu_result_6;
input 	r_sync_rst;
input 	d_write;
input 	write_accepted;
input 	rst1;
input 	cp_valid;
input 	F_pc_2;
input 	Equal4;
input 	cp_valid1;
output 	saved_grant_0;
output 	src_payload;
output 	saved_grant_1;
input 	Equal41;
output 	src_valid;
output 	src_valid1;
input 	uav_read;
input 	Equal42;
input 	uav_read1;
input 	src5_valid;
input 	write;
output 	WideOr11;
output 	src_data_56;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \src_valid~5_combout ;
wire \update_grant~0_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~1_combout ;
wire \src_valid~3_combout ;


processor_altera_merlin_arbitrator_4 arb(
	.reset(r_sync_rst),
	.src5_valid(src5_valid),
	.grant_0(\arb|grant[0]~0_combout ),
	.update_grant(\update_grant~1_combout ),
	.grant_1(\arb|grant[1]~1_combout ),
	.src_valid(\src_valid~5_combout ),
	.clk(clk_clk));

cyclone10lp_lcell_comb \src_valid~5 (
	.dataa(rst1),
	.datab(cp_valid1),
	.datac(Equal42),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_valid~5_combout ),
	.cout());
defparam \src_valid~5 .lut_mask = 16'hFBFB;
defparam \src_valid~5 .sum_lutc_input = "datac";

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

cyclone10lp_lcell_comb \src_payload~0 (
	.dataa(d_write),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(write_accepted),
	.cin(gnd),
	.combout(src_payload),
	.cout());
defparam \src_payload~0 .lut_mask = 16'hEEFF;
defparam \src_payload~0 .sum_lutc_input = "datac";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclone10lp_lcell_comb \src_valid~2 (
	.dataa(cp_valid),
	.datab(F_pc_2),
	.datac(saved_grant_1),
	.datad(Equal41),
	.cin(gnd),
	.combout(src_valid),
	.cout());
defparam \src_valid~2 .lut_mask = 16'hFFFE;
defparam \src_valid~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_valid~4 (
	.dataa(W_alu_result_4),
	.datab(Equal4),
	.datac(cp_valid1),
	.datad(\src_valid~3_combout ),
	.cin(gnd),
	.combout(src_valid1),
	.cout());
defparam \src_valid~4 .lut_mask = 16'hFFEF;
defparam \src_valid~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb WideOr1(
	.dataa(src_valid),
	.datab(src_valid1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam WideOr1.lut_mask = 16'hEEEE;
defparam WideOr1.sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[56] (
	.dataa(uav_read),
	.datab(uav_read1),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_56),
	.cout());
defparam \src_data[56] .lut_mask = 16'hFFFE;
defparam \src_data[56] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \update_grant~0 (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\update_grant~0_combout ),
	.cout());
defparam \update_grant~0 .lut_mask = 16'hEEEE;
defparam \update_grant~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \packet_in_progress~0 (
	.dataa(\update_grant~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\packet_in_progress~0_combout ),
	.cout());
defparam \packet_in_progress~0 .lut_mask = 16'h5555;
defparam \packet_in_progress~0 .sum_lutc_input = "datac";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclone10lp_lcell_comb \update_grant~1 (
	.dataa(\update_grant~0_combout ),
	.datab(write),
	.datac(WideOr11),
	.datad(\packet_in_progress~q ),
	.cin(gnd),
	.combout(\update_grant~1_combout ),
	.cout());
defparam \update_grant~1 .lut_mask = 16'hEFFF;
defparam \update_grant~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_valid~3 (
	.dataa(saved_grant_0),
	.datab(W_alu_result_5),
	.datac(W_alu_result_6),
	.datad(rst1),
	.cin(gnd),
	.combout(\src_valid~3_combout ),
	.cout());
defparam \src_valid~3 .lut_mask = 16'hFFBF;
defparam \src_valid~3 .sum_lutc_input = "datac";

endmodule

module processor_altera_merlin_arbitrator_4 (
	reset,
	src5_valid,
	grant_0,
	update_grant,
	grant_1,
	src_valid,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	src5_valid;
output 	grant_0;
input 	update_grant;
output 	grant_1;
input 	src_valid;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~q ;


cyclone10lp_lcell_comb \grant[0]~0 (
	.dataa(src_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(src5_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_0),
	.cout());
defparam \grant[0]~0 .lut_mask = 16'hEFFF;
defparam \grant[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \grant[1]~1 (
	.dataa(src5_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(src_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_1),
	.cout());
defparam \grant[1]~1 .lut_mask = 16'hEFFF;
defparam \grant[1]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \top_priority_reg[0]~0 (
	.dataa(update_grant),
	.datab(src5_valid),
	.datac(src_valid),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.cout());
defparam \top_priority_reg[0]~0 .lut_mask = 16'hFEFE;
defparam \top_priority_reg[0]~0 .sum_lutc_input = "datac";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cyclone10lp_lcell_comb \top_priority_reg[0]~1 (
	.dataa(grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.cout());
defparam \top_priority_reg[0]~1 .lut_mask = 16'h5555;
defparam \top_priority_reg[0]~1 .sum_lutc_input = "datac";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module processor_processor_mm_interconnect_0_cmd_mux_6 (
	W_alu_result_5,
	W_alu_result_6,
	r_sync_rst,
	rst1,
	cp_valid,
	Equal4,
	cp_valid1,
	Equal41,
	uav_read,
	always1,
	always11,
	saved_grant_0,
	always12,
	saved_grant_1,
	src_valid,
	src_valid1,
	always13,
	cp_ready,
	uav_read1,
	WideOr11,
	src_data_56,
	src6_valid,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_5;
input 	W_alu_result_6;
input 	r_sync_rst;
input 	rst1;
input 	cp_valid;
input 	Equal4;
input 	cp_valid1;
input 	Equal41;
input 	uav_read;
input 	always1;
input 	always11;
output 	saved_grant_0;
input 	always12;
output 	saved_grant_1;
output 	src_valid;
output 	src_valid1;
input 	always13;
input 	cp_ready;
input 	uav_read1;
output 	WideOr11;
output 	src_data_56;
input 	src6_valid;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \src_valid~5_combout ;
wire \update_grant~0_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~1_combout ;
wire \src_valid~3_combout ;


processor_altera_merlin_arbitrator_5 arb(
	.reset(r_sync_rst),
	.src6_valid(src6_valid),
	.grant_0(\arb|grant[0]~0_combout ),
	.update_grant(\update_grant~1_combout ),
	.grant_1(\arb|grant[1]~1_combout ),
	.src_valid(\src_valid~5_combout ),
	.clk(clk_clk));

cyclone10lp_lcell_comb \src_valid~5 (
	.dataa(rst1),
	.datab(cp_valid1),
	.datac(always11),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_valid~5_combout ),
	.cout());
defparam \src_valid~5 .lut_mask = 16'hFBFB;
defparam \src_valid~5 .sum_lutc_input = "datac";

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclone10lp_lcell_comb \src_valid~2 (
	.dataa(cp_valid),
	.datab(Equal41),
	.datac(always12),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_valid),
	.cout());
defparam \src_valid~2 .lut_mask = 16'hFFFE;
defparam \src_valid~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_valid~4 (
	.dataa(always1),
	.datab(Equal4),
	.datac(cp_valid1),
	.datad(\src_valid~3_combout ),
	.cin(gnd),
	.combout(src_valid1),
	.cout());
defparam \src_valid~4 .lut_mask = 16'hFFEF;
defparam \src_valid~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb WideOr1(
	.dataa(src_valid1),
	.datab(cp_valid),
	.datac(always13),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam WideOr1.lut_mask = 16'hFFFE;
defparam WideOr1.sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[56] (
	.dataa(uav_read),
	.datab(uav_read1),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_56),
	.cout());
defparam \src_data[56] .lut_mask = 16'hFFFE;
defparam \src_data[56] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \update_grant~0 (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\update_grant~0_combout ),
	.cout());
defparam \update_grant~0 .lut_mask = 16'hEEEE;
defparam \update_grant~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \packet_in_progress~0 (
	.dataa(\update_grant~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\packet_in_progress~0_combout ),
	.cout());
defparam \packet_in_progress~0 .lut_mask = 16'h5555;
defparam \packet_in_progress~0 .sum_lutc_input = "datac";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclone10lp_lcell_comb \update_grant~1 (
	.dataa(\update_grant~0_combout ),
	.datab(WideOr11),
	.datac(\packet_in_progress~q ),
	.datad(cp_ready),
	.cin(gnd),
	.combout(\update_grant~1_combout ),
	.cout());
defparam \update_grant~1 .lut_mask = 16'h8BFF;
defparam \update_grant~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_valid~3 (
	.dataa(saved_grant_0),
	.datab(W_alu_result_5),
	.datac(W_alu_result_6),
	.datad(rst1),
	.cin(gnd),
	.combout(\src_valid~3_combout ),
	.cout());
defparam \src_valid~3 .lut_mask = 16'hFFBF;
defparam \src_valid~3 .sum_lutc_input = "datac";

endmodule

module processor_altera_merlin_arbitrator_5 (
	reset,
	src6_valid,
	grant_0,
	update_grant,
	grant_1,
	src_valid,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	src6_valid;
output 	grant_0;
input 	update_grant;
output 	grant_1;
input 	src_valid;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~q ;


cyclone10lp_lcell_comb \grant[0]~0 (
	.dataa(src_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(src6_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_0),
	.cout());
defparam \grant[0]~0 .lut_mask = 16'hEFFF;
defparam \grant[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \grant[1]~1 (
	.dataa(src6_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(src_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_1),
	.cout());
defparam \grant[1]~1 .lut_mask = 16'hEFFF;
defparam \grant[1]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \top_priority_reg[0]~0 (
	.dataa(update_grant),
	.datab(src6_valid),
	.datac(src_valid),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.cout());
defparam \top_priority_reg[0]~0 .lut_mask = 16'hFEFE;
defparam \top_priority_reg[0]~0 .sum_lutc_input = "datac";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cyclone10lp_lcell_comb \top_priority_reg[0]~1 (
	.dataa(grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.cout());
defparam \top_priority_reg[0]~1 .lut_mask = 16'h5555;
defparam \top_priority_reg[0]~1 .sum_lutc_input = "datac";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module processor_processor_mm_interconnect_0_cmd_mux_7 (
	W_alu_result_4,
	W_alu_result_2,
	W_alu_result_3,
	d_writedata_0,
	r_sync_rst,
	rst1,
	F_pc_2,
	cp_valid,
	F_pc_1,
	F_pc_0,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	uav_read,
	Equal2,
	saved_grant_0,
	mem_used_1,
	uav_waitrequest,
	saved_grant_1,
	uav_read1,
	d_writedata_9,
	src_payload,
	src_data_38,
	src_data_39,
	src_data_40,
	WideOr11,
	src_data_56,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	d_writedata_8,
	src_payload9,
	src7_valid,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	W_alu_result_2;
input 	W_alu_result_3;
input 	d_writedata_0;
input 	r_sync_rst;
input 	rst1;
input 	F_pc_2;
input 	cp_valid;
input 	F_pc_1;
input 	F_pc_0;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
input 	uav_read;
input 	Equal2;
output 	saved_grant_0;
input 	mem_used_1;
input 	uav_waitrequest;
output 	saved_grant_1;
input 	uav_read1;
input 	d_writedata_9;
output 	src_payload;
output 	src_data_38;
output 	src_data_39;
output 	src_data_40;
output 	WideOr11;
output 	src_data_56;
output 	src_payload1;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
output 	src_payload7;
output 	src_payload8;
input 	d_writedata_8;
output 	src_payload9;
input 	src7_valid;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \update_grant~0_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~1_combout ;
wire \src_valid~2_combout ;


processor_altera_merlin_arbitrator_6 arb(
	.reset(r_sync_rst),
	.grant_0(\arb|grant[0]~0_combout ),
	.update_grant(\update_grant~1_combout ),
	.grant_1(\arb|grant[1]~1_combout ),
	.src_valid(\src_valid~2_combout ),
	.src7_valid(src7_valid),
	.clk(clk_clk));

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclone10lp_lcell_comb \src_payload~0 (
	.dataa(saved_grant_0),
	.datab(d_writedata_9),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload),
	.cout());
defparam \src_payload~0 .lut_mask = 16'hEEEE;
defparam \src_payload~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[38] (
	.dataa(W_alu_result_2),
	.datab(F_pc_0),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_38),
	.cout());
defparam \src_data[38] .lut_mask = 16'hFFFE;
defparam \src_data[38] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[39] (
	.dataa(W_alu_result_3),
	.datab(F_pc_1),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_39),
	.cout());
defparam \src_data[39] .lut_mask = 16'hFFFE;
defparam \src_data[39] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[40] (
	.dataa(F_pc_2),
	.datab(W_alu_result_4),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_40),
	.cout());
defparam \src_data[40] .lut_mask = 16'hFFFE;
defparam \src_data[40] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb WideOr1(
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(\src_valid~2_combout ),
	.datad(src7_valid),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam WideOr1.lut_mask = 16'hFFFE;
defparam WideOr1.sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[56] (
	.dataa(uav_read),
	.datab(uav_read1),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_56),
	.cout());
defparam \src_data[56] .lut_mask = 16'hFFFE;
defparam \src_data[56] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~1 (
	.dataa(d_writedata_7),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload1),
	.cout());
defparam \src_payload~1 .lut_mask = 16'hEEEE;
defparam \src_payload~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~2 (
	.dataa(d_writedata_6),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload2),
	.cout());
defparam \src_payload~2 .lut_mask = 16'hEEEE;
defparam \src_payload~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~3 (
	.dataa(d_writedata_5),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload3),
	.cout());
defparam \src_payload~3 .lut_mask = 16'hEEEE;
defparam \src_payload~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~4 (
	.dataa(d_writedata_4),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload4),
	.cout());
defparam \src_payload~4 .lut_mask = 16'hEEEE;
defparam \src_payload~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~5 (
	.dataa(d_writedata_3),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload5),
	.cout());
defparam \src_payload~5 .lut_mask = 16'hEEEE;
defparam \src_payload~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~6 (
	.dataa(d_writedata_2),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload6),
	.cout());
defparam \src_payload~6 .lut_mask = 16'hEEEE;
defparam \src_payload~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~7 (
	.dataa(d_writedata_1),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload7),
	.cout());
defparam \src_payload~7 .lut_mask = 16'hEEEE;
defparam \src_payload~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~8 (
	.dataa(d_writedata_0),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload8),
	.cout());
defparam \src_payload~8 .lut_mask = 16'hEEEE;
defparam \src_payload~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~9 (
	.dataa(saved_grant_0),
	.datab(d_writedata_8),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload9),
	.cout());
defparam \src_payload~9 .lut_mask = 16'hEEEE;
defparam \src_payload~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \update_grant~0 (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(uav_waitrequest),
	.cin(gnd),
	.combout(\update_grant~0_combout ),
	.cout());
defparam \update_grant~0 .lut_mask = 16'hEEFF;
defparam \update_grant~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \packet_in_progress~0 (
	.dataa(\update_grant~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\packet_in_progress~0_combout ),
	.cout());
defparam \packet_in_progress~0 .lut_mask = 16'h5555;
defparam \packet_in_progress~0 .sum_lutc_input = "datac";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclone10lp_lcell_comb \update_grant~1 (
	.dataa(\update_grant~0_combout ),
	.datab(WideOr11),
	.datac(\packet_in_progress~q ),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\update_grant~1_combout ),
	.cout());
defparam \update_grant~1 .lut_mask = 16'h8BFF;
defparam \update_grant~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_valid~2 (
	.dataa(rst1),
	.datab(cp_valid),
	.datac(Equal2),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_valid~2_combout ),
	.cout());
defparam \src_valid~2 .lut_mask = 16'hFBFB;
defparam \src_valid~2 .sum_lutc_input = "datac";

endmodule

module processor_altera_merlin_arbitrator_6 (
	reset,
	grant_0,
	update_grant,
	grant_1,
	src_valid,
	src7_valid,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
output 	grant_0;
input 	update_grant;
output 	grant_1;
input 	src_valid;
input 	src7_valid;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~q ;


cyclone10lp_lcell_comb \grant[0]~0 (
	.dataa(src_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(src7_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_0),
	.cout());
defparam \grant[0]~0 .lut_mask = 16'hEFFF;
defparam \grant[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \grant[1]~1 (
	.dataa(src7_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(src_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_1),
	.cout());
defparam \grant[1]~1 .lut_mask = 16'hEFFF;
defparam \grant[1]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \top_priority_reg[0]~0 (
	.dataa(update_grant),
	.datab(src7_valid),
	.datac(src_valid),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.cout());
defparam \top_priority_reg[0]~0 .lut_mask = 16'hFEFE;
defparam \top_priority_reg[0]~0 .sum_lutc_input = "datac";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cyclone10lp_lcell_comb \top_priority_reg[0]~1 (
	.dataa(grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.cout());
defparam \top_priority_reg[0]~1 .lut_mask = 16'h5555;
defparam \top_priority_reg[0]~1 .sum_lutc_input = "datac";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module processor_altera_merlin_arbitrator_7 (
	reset,
	src0_valid,
	grant_0,
	update_grant,
	grant_1,
	src_valid,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	src0_valid;
output 	grant_0;
input 	update_grant;
output 	grant_1;
input 	src_valid;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~q ;


cyclone10lp_lcell_comb \grant[0]~0 (
	.dataa(src_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(src0_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_0),
	.cout());
defparam \grant[0]~0 .lut_mask = 16'hEFFF;
defparam \grant[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \grant[1]~1 (
	.dataa(src0_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(src_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_1),
	.cout());
defparam \grant[1]~1 .lut_mask = 16'hEFFF;
defparam \grant[1]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \top_priority_reg[0]~0 (
	.dataa(update_grant),
	.datab(src0_valid),
	.datac(src_valid),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.cout());
defparam \top_priority_reg[0]~0 .lut_mask = 16'hFEFE;
defparam \top_priority_reg[0]~0 .sum_lutc_input = "datac";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cyclone10lp_lcell_comb \top_priority_reg[0]~1 (
	.dataa(grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.cout());
defparam \top_priority_reg[0]~1 .lut_mask = 16'h5555;
defparam \top_priority_reg[0]~1 .sum_lutc_input = "datac";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module processor_processor_mm_interconnect_0_router (
	W_alu_result_7,
	W_alu_result_16,
	W_alu_result_15,
	W_alu_result_14,
	W_alu_result_13,
	W_alu_result_12,
	W_alu_result_11,
	W_alu_result_10,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_4,
	W_alu_result_5,
	W_alu_result_6,
	W_alu_result_3,
	Equal4,
	read_accepted,
	d_read,
	Equal6,
	Equal5,
	Equal1,
	Equal7,
	Equal2,
	always1,
	always11,
	Equal41)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_7;
input 	W_alu_result_16;
input 	W_alu_result_15;
input 	W_alu_result_14;
input 	W_alu_result_13;
input 	W_alu_result_12;
input 	W_alu_result_11;
input 	W_alu_result_10;
input 	W_alu_result_9;
input 	W_alu_result_8;
input 	W_alu_result_4;
input 	W_alu_result_5;
input 	W_alu_result_6;
input 	W_alu_result_3;
output 	Equal4;
input 	read_accepted;
input 	d_read;
output 	Equal6;
output 	Equal5;
output 	Equal1;
output 	Equal7;
output 	Equal2;
output 	always1;
output 	always11;
output 	Equal41;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Equal1~0_combout ;
wire \Equal2~0_combout ;
wire \Equal6~0_combout ;
wire \Equal5~0_combout ;
wire \Equal2~1_combout ;


cyclone10lp_lcell_comb \Equal4~0 (
	.dataa(W_alu_result_7),
	.datab(\Equal1~0_combout ),
	.datac(\Equal2~0_combout ),
	.datad(W_alu_result_8),
	.cin(gnd),
	.combout(Equal4),
	.cout());
defparam \Equal4~0 .lut_mask = 16'hFEFF;
defparam \Equal4~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal6~1 (
	.dataa(W_alu_result_7),
	.datab(\Equal1~0_combout ),
	.datac(\Equal2~0_combout ),
	.datad(\Equal6~0_combout ),
	.cin(gnd),
	.combout(Equal6),
	.cout());
defparam \Equal6~1 .lut_mask = 16'hFFFE;
defparam \Equal6~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal5~1 (
	.dataa(W_alu_result_5),
	.datab(\Equal1~0_combout ),
	.datac(\Equal2~0_combout ),
	.datad(\Equal5~0_combout ),
	.cin(gnd),
	.combout(Equal5),
	.cout());
defparam \Equal5~1 .lut_mask = 16'hFFFE;
defparam \Equal5~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal1~1 (
	.dataa(W_alu_result_12),
	.datab(gnd),
	.datac(\Equal1~0_combout ),
	.datad(W_alu_result_11),
	.cin(gnd),
	.combout(Equal1),
	.cout());
defparam \Equal1~1 .lut_mask = 16'hAFFF;
defparam \Equal1~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal7~0 (
	.dataa(W_alu_result_6),
	.datab(W_alu_result_3),
	.datac(W_alu_result_4),
	.datad(W_alu_result_5),
	.cin(gnd),
	.combout(Equal7),
	.cout());
defparam \Equal7~0 .lut_mask = 16'hEFFF;
defparam \Equal7~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal2~2 (
	.dataa(\Equal1~0_combout ),
	.datab(\Equal2~0_combout ),
	.datac(\Equal2~1_combout ),
	.datad(W_alu_result_8),
	.cin(gnd),
	.combout(Equal2),
	.cout());
defparam \Equal2~2 .lut_mask = 16'hFEFF;
defparam \Equal2~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \always1~0 (
	.dataa(d_read),
	.datab(gnd),
	.datac(W_alu_result_4),
	.datad(read_accepted),
	.cin(gnd),
	.combout(always1),
	.cout());
defparam \always1~0 .lut_mask = 16'hAFFF;
defparam \always1~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \always1~1 (
	.dataa(Equal4),
	.datab(always1),
	.datac(W_alu_result_5),
	.datad(W_alu_result_6),
	.cin(gnd),
	.combout(always11),
	.cout());
defparam \always1~1 .lut_mask = 16'hEFFF;
defparam \always1~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal4~1 (
	.dataa(W_alu_result_4),
	.datab(Equal4),
	.datac(W_alu_result_5),
	.datad(W_alu_result_6),
	.cin(gnd),
	.combout(Equal41),
	.cout());
defparam \Equal4~1 .lut_mask = 16'hEFFF;
defparam \Equal4~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal1~0 (
	.dataa(W_alu_result_16),
	.datab(W_alu_result_15),
	.datac(W_alu_result_14),
	.datad(W_alu_result_13),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
defparam \Equal1~0 .lut_mask = 16'hBFFF;
defparam \Equal1~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal2~0 (
	.dataa(W_alu_result_12),
	.datab(W_alu_result_11),
	.datac(W_alu_result_10),
	.datad(W_alu_result_9),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
defparam \Equal2~0 .lut_mask = 16'hBFFF;
defparam \Equal2~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal6~0 (
	.dataa(W_alu_result_4),
	.datab(W_alu_result_5),
	.datac(W_alu_result_6),
	.datad(W_alu_result_8),
	.cin(gnd),
	.combout(\Equal6~0_combout ),
	.cout());
defparam \Equal6~0 .lut_mask = 16'hEFFF;
defparam \Equal6~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal5~0 (
	.dataa(W_alu_result_4),
	.datab(W_alu_result_6),
	.datac(W_alu_result_7),
	.datad(W_alu_result_8),
	.cin(gnd),
	.combout(\Equal5~0_combout ),
	.cout());
defparam \Equal5~0 .lut_mask = 16'hF7FF;
defparam \Equal5~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal2~1 (
	.dataa(W_alu_result_5),
	.datab(gnd),
	.datac(W_alu_result_6),
	.datad(W_alu_result_7),
	.cin(gnd),
	.combout(\Equal2~1_combout ),
	.cout());
defparam \Equal2~1 .lut_mask = 16'hAFFF;
defparam \Equal2~1 .sum_lutc_input = "datac";

endmodule

module processor_processor_mm_interconnect_0_router_1 (
	i_read,
	read_accepted,
	F_pc_5,
	F_pc_14,
	F_pc_13,
	F_pc_12,
	F_pc_11,
	Equal1,
	F_pc_10,
	F_pc_9,
	F_pc_8,
	F_pc_7,
	F_pc_6,
	Equal4,
	F_pc_2,
	F_pc_3,
	F_pc_4,
	F_pc_1,
	Equal41,
	Equal6,
	always1,
	Equal7,
	Equal11,
	src_channel_2,
	Equal2,
	src_channel_21,
	src_channel_22,
	Equal5,
	Equal42,
	always11)/* synthesis synthesis_greybox=1 */;
input 	i_read;
input 	read_accepted;
input 	F_pc_5;
input 	F_pc_14;
input 	F_pc_13;
input 	F_pc_12;
input 	F_pc_11;
output 	Equal1;
input 	F_pc_10;
input 	F_pc_9;
input 	F_pc_8;
input 	F_pc_7;
input 	F_pc_6;
output 	Equal4;
input 	F_pc_2;
input 	F_pc_3;
input 	F_pc_4;
input 	F_pc_1;
output 	Equal41;
output 	Equal6;
output 	always1;
output 	Equal7;
output 	Equal11;
output 	src_channel_2;
output 	Equal2;
output 	src_channel_21;
output 	src_channel_22;
output 	Equal5;
output 	Equal42;
output 	always11;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Equal2~0_combout ;
wire \Equal4~1_combout ;
wire \Equal6~0_combout ;
wire \Equal2~1_combout ;
wire \Equal5~0_combout ;


cyclone10lp_lcell_comb \Equal1~0 (
	.dataa(F_pc_14),
	.datab(F_pc_13),
	.datac(F_pc_12),
	.datad(F_pc_11),
	.cin(gnd),
	.combout(Equal1),
	.cout());
defparam \Equal1~0 .lut_mask = 16'hEFFF;
defparam \Equal1~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal4~0 (
	.dataa(F_pc_5),
	.datab(Equal1),
	.datac(\Equal2~0_combout ),
	.datad(F_pc_6),
	.cin(gnd),
	.combout(Equal4),
	.cout());
defparam \Equal4~0 .lut_mask = 16'hFEFF;
defparam \Equal4~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal4~2 (
	.dataa(F_pc_4),
	.datab(Equal1),
	.datac(\Equal2~0_combout ),
	.datad(\Equal4~1_combout ),
	.cin(gnd),
	.combout(Equal41),
	.cout());
defparam \Equal4~2 .lut_mask = 16'hFFFD;
defparam \Equal4~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal6~1 (
	.dataa(F_pc_5),
	.datab(Equal1),
	.datac(\Equal2~0_combout ),
	.datad(\Equal6~0_combout ),
	.cin(gnd),
	.combout(Equal6),
	.cout());
defparam \Equal6~1 .lut_mask = 16'hFFFE;
defparam \Equal6~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \always1~0 (
	.dataa(gnd),
	.datab(i_read),
	.datac(read_accepted),
	.datad(F_pc_2),
	.cin(gnd),
	.combout(always1),
	.cout());
defparam \always1~0 .lut_mask = 16'h3FFF;
defparam \always1~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal7~0 (
	.dataa(F_pc_4),
	.datab(F_pc_1),
	.datac(F_pc_2),
	.datad(F_pc_3),
	.cin(gnd),
	.combout(Equal7),
	.cout());
defparam \Equal7~0 .lut_mask = 16'hEFFF;
defparam \Equal7~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal1~1 (
	.dataa(F_pc_10),
	.datab(gnd),
	.datac(Equal1),
	.datad(F_pc_9),
	.cin(gnd),
	.combout(Equal11),
	.cout());
defparam \Equal1~1 .lut_mask = 16'hAFFF;
defparam \Equal1~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_channel[2]~0 (
	.dataa(F_pc_4),
	.datab(F_pc_2),
	.datac(F_pc_3),
	.datad(Equal4),
	.cin(gnd),
	.combout(src_channel_2),
	.cout());
defparam \src_channel[2]~0 .lut_mask = 16'hBFFF;
defparam \src_channel[2]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal2~2 (
	.dataa(Equal1),
	.datab(\Equal2~0_combout ),
	.datac(\Equal2~1_combout ),
	.datad(F_pc_6),
	.cin(gnd),
	.combout(Equal2),
	.cout());
defparam \Equal2~2 .lut_mask = 16'hFEFF;
defparam \Equal2~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_channel[2]~1 (
	.dataa(Equal11),
	.datab(Equal4),
	.datac(Equal7),
	.datad(Equal2),
	.cin(gnd),
	.combout(src_channel_21),
	.cout());
defparam \src_channel[2]~1 .lut_mask = 16'hBFFF;
defparam \src_channel[2]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_channel[2]~2 (
	.dataa(src_channel_2),
	.datab(src_channel_21),
	.datac(Equal41),
	.datad(always1),
	.cin(gnd),
	.combout(src_channel_22),
	.cout());
defparam \src_channel[2]~2 .lut_mask = 16'hEFFF;
defparam \src_channel[2]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal5~1 (
	.dataa(F_pc_3),
	.datab(Equal1),
	.datac(\Equal2~0_combout ),
	.datad(\Equal5~0_combout ),
	.cin(gnd),
	.combout(Equal5),
	.cout());
defparam \Equal5~1 .lut_mask = 16'hFFFE;
defparam \Equal5~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal4~3 (
	.dataa(F_pc_2),
	.datab(Equal4),
	.datac(F_pc_3),
	.datad(F_pc_4),
	.cin(gnd),
	.combout(Equal42),
	.cout());
defparam \Equal4~3 .lut_mask = 16'hEFFF;
defparam \Equal4~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \always1~1 (
	.dataa(Equal4),
	.datab(always1),
	.datac(F_pc_3),
	.datad(F_pc_4),
	.cin(gnd),
	.combout(always11),
	.cout());
defparam \always1~1 .lut_mask = 16'hEFFF;
defparam \always1~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal2~0 (
	.dataa(F_pc_10),
	.datab(F_pc_9),
	.datac(F_pc_8),
	.datad(F_pc_7),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
defparam \Equal2~0 .lut_mask = 16'hBFFF;
defparam \Equal2~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal4~1 (
	.dataa(F_pc_3),
	.datab(F_pc_5),
	.datac(F_pc_6),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal4~1_combout ),
	.cout());
defparam \Equal4~1 .lut_mask = 16'hDFDF;
defparam \Equal4~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal6~0 (
	.dataa(F_pc_2),
	.datab(F_pc_3),
	.datac(F_pc_4),
	.datad(F_pc_6),
	.cin(gnd),
	.combout(\Equal6~0_combout ),
	.cout());
defparam \Equal6~0 .lut_mask = 16'hEFFF;
defparam \Equal6~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal2~1 (
	.dataa(F_pc_3),
	.datab(gnd),
	.datac(F_pc_4),
	.datad(F_pc_5),
	.cin(gnd),
	.combout(\Equal2~1_combout ),
	.cout());
defparam \Equal2~1 .lut_mask = 16'hAFFF;
defparam \Equal2~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal5~0 (
	.dataa(F_pc_2),
	.datab(F_pc_4),
	.datac(F_pc_5),
	.datad(F_pc_6),
	.cin(gnd),
	.combout(\Equal5~0_combout ),
	.cout());
defparam \Equal5~0 .lut_mask = 16'hF7FF;
defparam \Equal5~0 .sum_lutc_input = "datac";

endmodule

module processor_processor_mm_interconnect_0_rsp_demux (
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	src0_valid,
	src1_valid)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	mem_74_0;
input 	mem_56_0;
output 	src0_valid;
output 	src1_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclone10lp_lcell_comb \src0_valid~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(gnd),
	.datac(mem_74_0),
	.datad(mem_56_0),
	.cin(gnd),
	.combout(src0_valid),
	.cout());
defparam \src0_valid~0 .lut_mask = 16'hAFFF;
defparam \src0_valid~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src1_valid~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(mem_74_0),
	.datac(mem_56_0),
	.datad(gnd),
	.cin(gnd),
	.combout(src1_valid),
	.cout());
defparam \src1_valid~0 .lut_mask = 16'hFEFE;
defparam \src1_valid~0 .sum_lutc_input = "datac";

endmodule

module processor_processor_mm_interconnect_0_rsp_demux_1 (
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	src0_valid,
	src1_valid)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	mem_74_0;
input 	mem_56_0;
output 	src0_valid;
output 	src1_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclone10lp_lcell_comb \src0_valid~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(gnd),
	.datac(mem_74_0),
	.datad(mem_56_0),
	.cin(gnd),
	.combout(src0_valid),
	.cout());
defparam \src0_valid~0 .lut_mask = 16'hAFFF;
defparam \src0_valid~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src1_valid~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(mem_74_0),
	.datac(mem_56_0),
	.datad(gnd),
	.cin(gnd),
	.combout(src1_valid),
	.cout());
defparam \src1_valid~0 .lut_mask = 16'hFEFE;
defparam \src1_valid~0 .sum_lutc_input = "datac";

endmodule

module processor_processor_mm_interconnect_0_rsp_demux_2 (
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	src0_valid,
	src1_valid)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	mem_74_0;
input 	mem_56_0;
output 	src0_valid;
output 	src1_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclone10lp_lcell_comb \src0_valid~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(gnd),
	.datac(mem_74_0),
	.datad(mem_56_0),
	.cin(gnd),
	.combout(src0_valid),
	.cout());
defparam \src0_valid~0 .lut_mask = 16'hAFFF;
defparam \src0_valid~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src1_valid~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(mem_74_0),
	.datac(mem_56_0),
	.datad(gnd),
	.cin(gnd),
	.combout(src1_valid),
	.cout());
defparam \src1_valid~0 .lut_mask = 16'hFEFE;
defparam \src1_valid~0 .sum_lutc_input = "datac";

endmodule

module processor_processor_mm_interconnect_0_rsp_demux_3 (
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	src0_valid)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	mem_74_0;
input 	mem_56_0;
output 	src0_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclone10lp_lcell_comb \src0_valid~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(gnd),
	.datac(mem_74_0),
	.datad(mem_56_0),
	.cin(gnd),
	.combout(src0_valid),
	.cout());
defparam \src0_valid~0 .lut_mask = 16'hAFFF;
defparam \src0_valid~0 .sum_lutc_input = "datac";

endmodule

module processor_processor_mm_interconnect_0_rsp_demux_4 (
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	src0_valid)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	mem_74_0;
input 	mem_56_0;
output 	src0_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclone10lp_lcell_comb \src0_valid~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(gnd),
	.datac(mem_74_0),
	.datad(mem_56_0),
	.cin(gnd),
	.combout(src0_valid),
	.cout());
defparam \src0_valid~0 .lut_mask = 16'hAFFF;
defparam \src0_valid~0 .sum_lutc_input = "datac";

endmodule

module processor_processor_mm_interconnect_0_rsp_demux_5 (
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	src0_valid,
	src1_valid)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	mem_74_0;
input 	mem_56_0;
output 	src0_valid;
output 	src1_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclone10lp_lcell_comb \src0_valid~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(gnd),
	.datac(mem_74_0),
	.datad(mem_56_0),
	.cin(gnd),
	.combout(src0_valid),
	.cout());
defparam \src0_valid~0 .lut_mask = 16'hAFFF;
defparam \src0_valid~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src1_valid~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(mem_74_0),
	.datac(mem_56_0),
	.datad(gnd),
	.cin(gnd),
	.combout(src1_valid),
	.cout());
defparam \src1_valid~0 .lut_mask = 16'hFEFE;
defparam \src1_valid~0 .sum_lutc_input = "datac";

endmodule

module processor_processor_mm_interconnect_0_rsp_demux_6 (
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	src0_valid)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	mem_74_0;
input 	mem_56_0;
output 	src0_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclone10lp_lcell_comb \src0_valid~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(gnd),
	.datac(mem_74_0),
	.datad(mem_56_0),
	.cin(gnd),
	.combout(src0_valid),
	.cout());
defparam \src0_valid~0 .lut_mask = 16'hAFFF;
defparam \src0_valid~0 .sum_lutc_input = "datac";

endmodule

module processor_processor_mm_interconnect_0_rsp_demux_7 (
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	src0_valid,
	src1_valid)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	mem_74_0;
input 	mem_56_0;
output 	src0_valid;
output 	src1_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclone10lp_lcell_comb \src0_valid~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(gnd),
	.datac(mem_74_0),
	.datad(mem_56_0),
	.cin(gnd),
	.combout(src0_valid),
	.cout());
defparam \src0_valid~0 .lut_mask = 16'hAFFF;
defparam \src0_valid~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src1_valid~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(mem_74_0),
	.datac(mem_56_0),
	.datad(gnd),
	.cin(gnd),
	.combout(src1_valid),
	.cout());
defparam \src1_valid~0 .lut_mask = 16'hFEFE;
defparam \src1_valid~0 .sum_lutc_input = "datac";

endmodule

module processor_processor_mm_interconnect_0_rsp_mux (
	q_a_0,
	q_a_22,
	av_readdata_pre_22,
	q_a_23,
	q_a_14,
	q_a_15,
	q_a_11,
	q_a_13,
	q_a_16,
	av_readdata_pre_16,
	q_a_12,
	q_a_10,
	q_a_9,
	q_a_8,
	q_a_21,
	av_readdata_pre_21,
	q_a_20,
	av_readdata_pre_20,
	q_a_19,
	av_readdata_pre_19,
	q_a_18,
	av_readdata_pre_18,
	q_a_17,
	av_readdata_pre_17,
	src0_valid,
	src0_valid1,
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	src0_valid2,
	src0_valid3,
	WideOr11,
	src0_valid4,
	src0_valid5,
	src0_valid6,
	src0_valid7,
	WideOr12,
	WideOr13,
	av_readdata_pre_0,
	av_readdata_pre_01,
	av_readdata_pre_02,
	av_readdata_pre_03,
	av_readdata_pre_04,
	av_readdata_pre_05,
	av_readdata_pre_06,
	src_data_0,
	av_readdata_pre_221,
	av_readdata_pre_23,
	av_readdata_pre_14,
	av_readdata_pre_141,
	av_readdata_pre_15,
	av_readdata_pre_151,
	av_readdata_pre_11,
	av_readdata_pre_13,
	av_readdata_pre_131,
	av_readdata_pre_161,
	av_readdata_pre_12,
	av_readdata_pre_121,
	av_readdata_pre_10,
	av_readdata_pre_101,
	av_readdata_pre_9,
	av_readdata_pre_91,
	av_readdata_pre_92,
	av_readdata_pre_8,
	av_readdata_pre_81,
	av_readdata_pre_82,
	av_readdata_pre_211,
	av_readdata_pre_201,
	av_readdata_pre_191,
	av_readdata_pre_181,
	av_readdata_pre_171,
	src_data_8,
	src_payload,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_data_9,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13)/* synthesis synthesis_greybox=1 */;
input 	q_a_0;
input 	q_a_22;
input 	av_readdata_pre_22;
input 	q_a_23;
input 	q_a_14;
input 	q_a_15;
input 	q_a_11;
input 	q_a_13;
input 	q_a_16;
input 	av_readdata_pre_16;
input 	q_a_12;
input 	q_a_10;
input 	q_a_9;
input 	q_a_8;
input 	q_a_21;
input 	av_readdata_pre_21;
input 	q_a_20;
input 	av_readdata_pre_20;
input 	q_a_19;
input 	av_readdata_pre_19;
input 	q_a_18;
input 	av_readdata_pre_18;
input 	q_a_17;
input 	av_readdata_pre_17;
input 	src0_valid;
input 	src0_valid1;
input 	read_latency_shift_reg_0;
input 	mem_74_0;
input 	mem_56_0;
input 	src0_valid2;
input 	src0_valid3;
output 	WideOr11;
input 	src0_valid4;
input 	src0_valid5;
input 	src0_valid6;
input 	src0_valid7;
output 	WideOr12;
output 	WideOr13;
input 	av_readdata_pre_0;
input 	av_readdata_pre_01;
input 	av_readdata_pre_02;
input 	av_readdata_pre_03;
input 	av_readdata_pre_04;
input 	av_readdata_pre_05;
input 	av_readdata_pre_06;
output 	src_data_0;
input 	av_readdata_pre_221;
input 	av_readdata_pre_23;
input 	av_readdata_pre_14;
input 	av_readdata_pre_141;
input 	av_readdata_pre_15;
input 	av_readdata_pre_151;
input 	av_readdata_pre_11;
input 	av_readdata_pre_13;
input 	av_readdata_pre_131;
input 	av_readdata_pre_161;
input 	av_readdata_pre_12;
input 	av_readdata_pre_121;
input 	av_readdata_pre_10;
input 	av_readdata_pre_101;
input 	av_readdata_pre_9;
input 	av_readdata_pre_91;
input 	av_readdata_pre_92;
input 	av_readdata_pre_8;
input 	av_readdata_pre_81;
input 	av_readdata_pre_82;
input 	av_readdata_pre_211;
input 	av_readdata_pre_201;
input 	av_readdata_pre_191;
input 	av_readdata_pre_181;
input 	av_readdata_pre_171;
output 	src_data_8;
output 	src_payload;
output 	src_payload1;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
output 	src_data_9;
output 	src_payload7;
output 	src_payload8;
output 	src_payload9;
output 	src_payload10;
output 	src_payload11;
output 	src_payload12;
output 	src_payload13;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \src_data[0]~0_combout ;
wire \src_data[0]~1_combout ;
wire \src_data[0]~2_combout ;
wire \src_data[0]~3_combout ;
wire \src_data[8]~4_combout ;
wire \src_payload~0_combout ;
wire \src_payload~1_combout ;
wire \src_payload~3_combout ;
wire \src_payload~5_combout ;
wire \src_payload~7_combout ;
wire \src_payload~9_combout ;
wire \src_payload~12_combout ;
wire \src_data[9]~6_combout ;
wire \src_data[9]~7_combout ;
wire \src_payload~15_combout ;
wire \src_payload~17_combout ;
wire \src_payload~19_combout ;
wire \src_payload~21_combout ;
wire \src_payload~23_combout ;
wire \src_payload~25_combout ;


cyclone10lp_lcell_comb \WideOr1~0 (
	.dataa(src0_valid),
	.datab(src0_valid1),
	.datac(src0_valid2),
	.datad(src0_valid3),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam \WideOr1~0 .lut_mask = 16'h7FFF;
defparam \WideOr1~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \WideOr1~1 (
	.dataa(src0_valid4),
	.datab(src0_valid5),
	.datac(src0_valid6),
	.datad(src0_valid7),
	.cin(gnd),
	.combout(WideOr12),
	.cout());
defparam \WideOr1~1 .lut_mask = 16'h7FFF;
defparam \WideOr1~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb WideOr1(
	.dataa(WideOr11),
	.datab(WideOr12),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(WideOr13),
	.cout());
defparam WideOr1.lut_mask = 16'hEEEE;
defparam WideOr1.sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[0] (
	.dataa(\src_data[0]~0_combout ),
	.datab(src0_valid2),
	.datac(q_a_0),
	.datad(\src_data[0]~3_combout ),
	.cin(gnd),
	.combout(src_data_0),
	.cout());
defparam \src_data[0] .lut_mask = 16'hFFFE;
defparam \src_data[0] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[8]~5 (
	.dataa(\src_data[8]~4_combout ),
	.datab(\src_payload~0_combout ),
	.datac(src0_valid7),
	.datad(av_readdata_pre_82),
	.cin(gnd),
	.combout(src_data_8),
	.cout());
defparam \src_data[8]~5 .lut_mask = 16'hFFFE;
defparam \src_data[8]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~2 (
	.dataa(src0_valid2),
	.datab(q_a_16),
	.datac(\src_payload~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload),
	.cout());
defparam \src_payload~2 .lut_mask = 16'hFEFE;
defparam \src_payload~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~4 (
	.dataa(src0_valid2),
	.datab(q_a_15),
	.datac(\src_payload~3_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload1),
	.cout());
defparam \src_payload~4 .lut_mask = 16'hFEFE;
defparam \src_payload~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~6 (
	.dataa(src0_valid2),
	.datab(q_a_14),
	.datac(\src_payload~5_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload2),
	.cout());
defparam \src_payload~6 .lut_mask = 16'hFEFE;
defparam \src_payload~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~8 (
	.dataa(src0_valid2),
	.datab(q_a_13),
	.datac(\src_payload~7_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload3),
	.cout());
defparam \src_payload~8 .lut_mask = 16'hFEFE;
defparam \src_payload~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~10 (
	.dataa(src0_valid2),
	.datab(q_a_12),
	.datac(\src_payload~9_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload4),
	.cout());
defparam \src_payload~10 .lut_mask = 16'hFEFE;
defparam \src_payload~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~11 (
	.dataa(src0_valid1),
	.datab(src0_valid2),
	.datac(q_a_11),
	.datad(av_readdata_pre_11),
	.cin(gnd),
	.combout(src_payload5),
	.cout());
defparam \src_payload~11 .lut_mask = 16'hFFFE;
defparam \src_payload~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~13 (
	.dataa(src0_valid2),
	.datab(q_a_10),
	.datac(\src_payload~12_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload6),
	.cout());
defparam \src_payload~13 .lut_mask = 16'hFEFE;
defparam \src_payload~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[9]~8 (
	.dataa(src0_valid),
	.datab(av_readdata_pre_91),
	.datac(\src_data[9]~6_combout ),
	.datad(\src_data[9]~7_combout ),
	.cin(gnd),
	.combout(src_data_9),
	.cout());
defparam \src_data[9]~8 .lut_mask = 16'hFFFE;
defparam \src_data[9]~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~14 (
	.dataa(src0_valid1),
	.datab(src0_valid2),
	.datac(q_a_23),
	.datad(av_readdata_pre_23),
	.cin(gnd),
	.combout(src_payload7),
	.cout());
defparam \src_payload~14 .lut_mask = 16'hFFFE;
defparam \src_payload~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~16 (
	.dataa(src0_valid2),
	.datab(q_a_22),
	.datac(\src_payload~15_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload8),
	.cout());
defparam \src_payload~16 .lut_mask = 16'hFEFE;
defparam \src_payload~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~18 (
	.dataa(src0_valid2),
	.datab(q_a_21),
	.datac(\src_payload~17_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload9),
	.cout());
defparam \src_payload~18 .lut_mask = 16'hFEFE;
defparam \src_payload~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~20 (
	.dataa(src0_valid2),
	.datab(q_a_20),
	.datac(\src_payload~19_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload10),
	.cout());
defparam \src_payload~20 .lut_mask = 16'hFEFE;
defparam \src_payload~20 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~22 (
	.dataa(src0_valid2),
	.datab(q_a_19),
	.datac(\src_payload~21_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload11),
	.cout());
defparam \src_payload~22 .lut_mask = 16'hFEFE;
defparam \src_payload~22 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~24 (
	.dataa(src0_valid2),
	.datab(q_a_18),
	.datac(\src_payload~23_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload12),
	.cout());
defparam \src_payload~24 .lut_mask = 16'hFEFE;
defparam \src_payload~24 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~26 (
	.dataa(src0_valid2),
	.datab(q_a_17),
	.datac(\src_payload~25_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload13),
	.cout());
defparam \src_payload~26 .lut_mask = 16'hFEFE;
defparam \src_payload~26 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[0]~0 (
	.dataa(src0_valid4),
	.datab(src0_valid5),
	.datac(av_readdata_pre_0),
	.datad(av_readdata_pre_01),
	.cin(gnd),
	.combout(\src_data[0]~0_combout ),
	.cout());
defparam \src_data[0]~0 .lut_mask = 16'hFFFE;
defparam \src_data[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[0]~1 (
	.dataa(src0_valid1),
	.datab(av_readdata_pre_03),
	.datac(src0_valid7),
	.datad(av_readdata_pre_04),
	.cin(gnd),
	.combout(\src_data[0]~1_combout ),
	.cout());
defparam \src_data[0]~1 .lut_mask = 16'hFFFE;
defparam \src_data[0]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[0]~2 (
	.dataa(src0_valid3),
	.datab(av_readdata_pre_05),
	.datac(src0_valid6),
	.datad(av_readdata_pre_06),
	.cin(gnd),
	.combout(\src_data[0]~2_combout ),
	.cout());
defparam \src_data[0]~2 .lut_mask = 16'hFFFE;
defparam \src_data[0]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[0]~3 (
	.dataa(src0_valid),
	.datab(av_readdata_pre_02),
	.datac(\src_data[0]~1_combout ),
	.datad(\src_data[0]~2_combout ),
	.cin(gnd),
	.combout(\src_data[0]~3_combout ),
	.cout());
defparam \src_data[0]~3 .lut_mask = 16'hFFFE;
defparam \src_data[0]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[8]~4 (
	.dataa(src0_valid),
	.datab(src0_valid1),
	.datac(av_readdata_pre_8),
	.datad(av_readdata_pre_81),
	.cin(gnd),
	.combout(\src_data[8]~4_combout ),
	.cout());
defparam \src_data[8]~4 .lut_mask = 16'hFFFE;
defparam \src_data[8]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(q_a_8),
	.datac(mem_74_0),
	.datad(mem_56_0),
	.cin(gnd),
	.combout(\src_payload~0_combout ),
	.cout());
defparam \src_payload~0 .lut_mask = 16'hEFFF;
defparam \src_payload~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~1 (
	.dataa(src0_valid),
	.datab(av_readdata_pre_16),
	.datac(src0_valid1),
	.datad(av_readdata_pre_161),
	.cin(gnd),
	.combout(\src_payload~1_combout ),
	.cout());
defparam \src_payload~1 .lut_mask = 16'hFFFE;
defparam \src_payload~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~3 (
	.dataa(src0_valid),
	.datab(av_readdata_pre_151),
	.datac(src0_valid1),
	.datad(av_readdata_pre_15),
	.cin(gnd),
	.combout(\src_payload~3_combout ),
	.cout());
defparam \src_payload~3 .lut_mask = 16'hFFFE;
defparam \src_payload~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~5 (
	.dataa(src0_valid),
	.datab(av_readdata_pre_141),
	.datac(src0_valid1),
	.datad(av_readdata_pre_14),
	.cin(gnd),
	.combout(\src_payload~5_combout ),
	.cout());
defparam \src_payload~5 .lut_mask = 16'hFFFE;
defparam \src_payload~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~7 (
	.dataa(src0_valid),
	.datab(av_readdata_pre_131),
	.datac(src0_valid1),
	.datad(av_readdata_pre_13),
	.cin(gnd),
	.combout(\src_payload~7_combout ),
	.cout());
defparam \src_payload~7 .lut_mask = 16'hFFFE;
defparam \src_payload~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~9 (
	.dataa(src0_valid),
	.datab(av_readdata_pre_121),
	.datac(src0_valid1),
	.datad(av_readdata_pre_12),
	.cin(gnd),
	.combout(\src_payload~9_combout ),
	.cout());
defparam \src_payload~9 .lut_mask = 16'hFFFE;
defparam \src_payload~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~12 (
	.dataa(src0_valid),
	.datab(av_readdata_pre_101),
	.datac(src0_valid1),
	.datad(av_readdata_pre_10),
	.cin(gnd),
	.combout(\src_payload~12_combout ),
	.cout());
defparam \src_payload~12 .lut_mask = 16'hFFFE;
defparam \src_payload~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[9]~6 (
	.dataa(src0_valid7),
	.datab(av_readdata_pre_92),
	.datac(src0_valid1),
	.datad(av_readdata_pre_9),
	.cin(gnd),
	.combout(\src_data[9]~6_combout ),
	.cout());
defparam \src_data[9]~6 .lut_mask = 16'hFFFE;
defparam \src_data[9]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[9]~7 (
	.dataa(mem_74_0),
	.datab(mem_56_0),
	.datac(read_latency_shift_reg_0),
	.datad(q_a_9),
	.cin(gnd),
	.combout(\src_data[9]~7_combout ),
	.cout());
defparam \src_data[9]~7 .lut_mask = 16'hFFF7;
defparam \src_data[9]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~15 (
	.dataa(src0_valid),
	.datab(av_readdata_pre_22),
	.datac(src0_valid1),
	.datad(av_readdata_pre_221),
	.cin(gnd),
	.combout(\src_payload~15_combout ),
	.cout());
defparam \src_payload~15 .lut_mask = 16'hFFFE;
defparam \src_payload~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~17 (
	.dataa(src0_valid),
	.datab(av_readdata_pre_21),
	.datac(src0_valid1),
	.datad(av_readdata_pre_211),
	.cin(gnd),
	.combout(\src_payload~17_combout ),
	.cout());
defparam \src_payload~17 .lut_mask = 16'hFFFE;
defparam \src_payload~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~19 (
	.dataa(src0_valid),
	.datab(av_readdata_pre_20),
	.datac(src0_valid1),
	.datad(av_readdata_pre_201),
	.cin(gnd),
	.combout(\src_payload~19_combout ),
	.cout());
defparam \src_payload~19 .lut_mask = 16'hFFFE;
defparam \src_payload~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~21 (
	.dataa(src0_valid),
	.datab(av_readdata_pre_19),
	.datac(src0_valid1),
	.datad(av_readdata_pre_191),
	.cin(gnd),
	.combout(\src_payload~21_combout ),
	.cout());
defparam \src_payload~21 .lut_mask = 16'hFFFE;
defparam \src_payload~21 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~23 (
	.dataa(src0_valid),
	.datab(av_readdata_pre_18),
	.datac(src0_valid1),
	.datad(av_readdata_pre_181),
	.cin(gnd),
	.combout(\src_payload~23_combout ),
	.cout());
defparam \src_payload~23 .lut_mask = 16'hFFFE;
defparam \src_payload~23 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~25 (
	.dataa(src0_valid),
	.datab(av_readdata_pre_17),
	.datac(src0_valid1),
	.datad(av_readdata_pre_171),
	.cin(gnd),
	.combout(\src_payload~25_combout ),
	.cout());
defparam \src_payload~25 .lut_mask = 16'hFFFE;
defparam \src_payload~25 .sum_lutc_input = "datac";

endmodule

module processor_processor_mm_interconnect_0_rsp_mux_1 (
	q_a_0,
	q_a_11,
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	read_latency_shift_reg_01,
	mem_74_01,
	mem_56_01,
	read_latency_shift_reg_02,
	mem_74_02,
	mem_56_02,
	read_latency_shift_reg_03,
	mem_74_03,
	mem_56_03,
	read_latency_shift_reg_04,
	mem_74_04,
	mem_56_04,
	src1_valid,
	src1_valid1,
	src1_valid2,
	src1_valid3,
	WideOr1,
	src1_valid4,
	src_payload,
	src_payload1,
	WideOr11,
	av_readdata_pre_0,
	av_readdata_pre_01,
	av_readdata_pre_02,
	av_readdata_pre_03,
	av_readdata_pre_04,
	av_readdata_pre_05,
	av_readdata_pre_06,
	src_data_0,
	src_data_01,
	src_data_02,
	av_readdata_pre_3,
	src_payload2,
	src_payload3)/* synthesis synthesis_greybox=1 */;
input 	q_a_0;
input 	q_a_11;
input 	read_latency_shift_reg_0;
input 	mem_74_0;
input 	mem_56_0;
input 	read_latency_shift_reg_01;
input 	mem_74_01;
input 	mem_56_01;
input 	read_latency_shift_reg_02;
input 	mem_74_02;
input 	mem_56_02;
input 	read_latency_shift_reg_03;
input 	mem_74_03;
input 	mem_56_03;
input 	read_latency_shift_reg_04;
input 	mem_74_04;
input 	mem_56_04;
input 	src1_valid;
input 	src1_valid1;
input 	src1_valid2;
input 	src1_valid3;
output 	WideOr1;
input 	src1_valid4;
output 	src_payload;
output 	src_payload1;
output 	WideOr11;
input 	av_readdata_pre_0;
input 	av_readdata_pre_01;
input 	av_readdata_pre_02;
input 	av_readdata_pre_03;
input 	av_readdata_pre_04;
input 	av_readdata_pre_05;
input 	av_readdata_pre_06;
output 	src_data_0;
output 	src_data_01;
output 	src_data_02;
input 	av_readdata_pre_3;
output 	src_payload2;
output 	src_payload3;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \src_payload~2_combout ;
wire \src_data[0]~2_combout ;
wire \src_payload~3_combout ;


cyclone10lp_lcell_comb \WideOr1~0 (
	.dataa(src1_valid),
	.datab(src1_valid1),
	.datac(src1_valid2),
	.datad(src1_valid3),
	.cin(gnd),
	.combout(WideOr1),
	.cout());
defparam \WideOr1~0 .lut_mask = 16'hFFFE;
defparam \WideOr1~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~0 (
	.dataa(read_latency_shift_reg_03),
	.datab(mem_74_03),
	.datac(mem_56_03),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload),
	.cout());
defparam \src_payload~0 .lut_mask = 16'hFEFE;
defparam \src_payload~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~1 (
	.dataa(read_latency_shift_reg_02),
	.datab(mem_74_02),
	.datac(mem_56_02),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload1),
	.cout());
defparam \src_payload~1 .lut_mask = 16'hFEFE;
defparam \src_payload~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \WideOr1~1 (
	.dataa(src1_valid4),
	.datab(src_payload),
	.datac(src_payload1),
	.datad(\src_payload~2_combout ),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam \WideOr1~1 .lut_mask = 16'hFFFE;
defparam \WideOr1~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[0]~0 (
	.dataa(src1_valid),
	.datab(src1_valid1),
	.datac(av_readdata_pre_03),
	.datad(av_readdata_pre_02),
	.cin(gnd),
	.combout(src_data_0),
	.cout());
defparam \src_data[0]~0 .lut_mask = 16'hFFFE;
defparam \src_data[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[0]~1 (
	.dataa(src1_valid2),
	.datab(src1_valid3),
	.datac(av_readdata_pre_0),
	.datad(q_a_0),
	.cin(gnd),
	.combout(src_data_01),
	.cout());
defparam \src_data[0]~1 .lut_mask = 16'hFFFE;
defparam \src_data[0]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[0]~3 (
	.dataa(\src_data[0]~2_combout ),
	.datab(\src_payload~3_combout ),
	.datac(src_payload),
	.datad(av_readdata_pre_01),
	.cin(gnd),
	.combout(src_data_02),
	.cout());
defparam \src_data[0]~3 .lut_mask = 16'hFFFE;
defparam \src_data[0]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~4 (
	.dataa(read_latency_shift_reg_0),
	.datab(mem_74_0),
	.datac(mem_56_0),
	.datad(av_readdata_pre_3),
	.cin(gnd),
	.combout(src_payload2),
	.cout());
defparam \src_payload~4 .lut_mask = 16'hFFFE;
defparam \src_payload~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~5 (
	.dataa(read_latency_shift_reg_01),
	.datab(mem_74_01),
	.datac(mem_56_01),
	.datad(q_a_11),
	.cin(gnd),
	.combout(src_payload3),
	.cout());
defparam \src_payload~5 .lut_mask = 16'hFFFE;
defparam \src_payload~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~2 (
	.dataa(read_latency_shift_reg_04),
	.datab(mem_74_04),
	.datac(mem_56_04),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_payload~2_combout ),
	.cout());
defparam \src_payload~2 .lut_mask = 16'hFEFE;
defparam \src_payload~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_data[0]~2 (
	.dataa(src1_valid4),
	.datab(src_payload1),
	.datac(av_readdata_pre_05),
	.datad(av_readdata_pre_04),
	.cin(gnd),
	.combout(\src_data[0]~2_combout ),
	.cout());
defparam \src_data[0]~2 .lut_mask = 16'hFFFE;
defparam \src_data[0]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \src_payload~3 (
	.dataa(read_latency_shift_reg_04),
	.datab(mem_74_04),
	.datac(mem_56_04),
	.datad(av_readdata_pre_06),
	.cin(gnd),
	.combout(\src_payload~3_combout ),
	.cout());
defparam \src_payload~3 .lut_mask = 16'hFFFE;
defparam \src_payload~3 .sum_lutc_input = "datac";

endmodule

module processor_processor_nios2_gen2_0 (
	sr_0,
	W_alu_result_7,
	W_alu_result_16,
	W_alu_result_15,
	W_alu_result_14,
	W_alu_result_13,
	W_alu_result_12,
	W_alu_result_11,
	W_alu_result_10,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_4,
	W_alu_result_5,
	W_alu_result_6,
	W_alu_result_2,
	W_alu_result_3,
	q_a_22,
	av_readdata_pre_22,
	q_a_23,
	q_a_24,
	q_a_25,
	q_a_26,
	q_a_1,
	q_a_4,
	q_a_3,
	q_a_2,
	q_a_5,
	q_a_14,
	q_a_15,
	q_a_13,
	q_a_16,
	av_readdata_pre_16,
	q_a_12,
	q_a_10,
	q_a_9,
	q_a_8,
	q_a_7,
	q_a_6,
	q_a_21,
	av_readdata_pre_21,
	q_a_20,
	av_readdata_pre_20,
	q_a_19,
	av_readdata_pre_19,
	q_a_18,
	av_readdata_pre_18,
	q_a_17,
	av_readdata_pre_17,
	readdata_0,
	d_writedata_24,
	d_writedata_25,
	d_writedata_26,
	readdata_1,
	readdata_3,
	readdata_2,
	q_a_27,
	q_a_28,
	q_a_29,
	q_a_30,
	q_a_31,
	d_writedata_27,
	d_writedata_28,
	d_writedata_29,
	d_writedata_30,
	d_writedata_31,
	ir_out_0,
	ir_out_1,
	d_writedata_0,
	r_sync_rst,
	d_write,
	i_read,
	F_pc_5,
	F_pc_14,
	F_pc_13,
	F_pc_12,
	F_pc_11,
	F_pc_10,
	F_pc_9,
	F_pc_8,
	F_pc_7,
	F_pc_6,
	F_pc_2,
	F_pc_3,
	F_pc_4,
	d_read,
	F_pc_1,
	F_pc_0,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	src0_valid,
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	src0_valid1,
	read_latency_shift_reg_01,
	mem_74_01,
	mem_56_01,
	src0_valid2,
	src0_valid3,
	WideOr1,
	src0_valid4,
	read_latency_shift_reg_02,
	mem_74_02,
	mem_56_02,
	src0_valid5,
	src0_valid6,
	WideOr11,
	WideOr12,
	saved_grant_0,
	debug_mem_slave_waitrequest,
	mem_used_1,
	av_waitrequest,
	src1_valid,
	src1_valid1,
	src1_valid2,
	src1_valid3,
	WideOr13,
	src1_valid4,
	src_payload,
	src_payload1,
	WideOr14,
	uav_write,
	d_writedata_9,
	WideOr15,
	rf_source_valid,
	hbreak_enabled,
	src_data_0,
	av_readdata_pre_221,
	av_readdata_pre_23,
	av_readdata_pre_24,
	av_readdata_pre_25,
	av_readdata_pre_26,
	src_data_01,
	src_data_02,
	src_data_03,
	av_readdata_pre_1,
	av_readdata_pre_11,
	av_readdata_pre_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	av_readdata_pre_15,
	av_readdata_pre_4,
	av_readdata_pre_41,
	av_readdata_pre_42,
	av_readdata_pre_43,
	av_readdata_pre_3,
	src_payload2,
	av_readdata_pre_31,
	av_readdata_pre_32,
	av_readdata_pre_33,
	av_readdata_pre_2,
	av_readdata_pre_27,
	av_readdata_pre_28,
	av_readdata_pre_29,
	av_readdata_pre_210,
	src_data_46,
	av_readdata_pre_5,
	av_readdata_pre_51,
	av_readdata_pre_52,
	av_readdata_pre_53,
	av_readdata_pre_141,
	av_readdata_pre_142,
	av_readdata_pre_151,
	av_readdata_pre_152,
	src_payload3,
	av_readdata_pre_111,
	av_readdata_pre_131,
	av_readdata_pre_132,
	av_readdata_pre_161,
	av_readdata_pre_121,
	av_readdata_pre_122,
	av_readdata_pre_10,
	av_readdata_pre_101,
	av_readdata_pre_9,
	av_readdata_pre_91,
	av_readdata_pre_92,
	av_readdata_pre_8,
	av_readdata_pre_81,
	av_readdata_pre_82,
	av_readdata_pre_7,
	av_readdata_pre_71,
	av_readdata_pre_72,
	av_readdata_pre_73,
	av_readdata_pre_6,
	av_readdata_pre_61,
	av_readdata_pre_62,
	av_readdata_pre_63,
	av_readdata_pre_211,
	av_readdata_pre_201,
	av_readdata_pre_191,
	av_readdata_pre_181,
	av_readdata_pre_171,
	r_early_rst,
	src_data_8,
	d_byteenable_0,
	av_readdata_9,
	av_readdata_8,
	irq,
	d_writedata_22,
	d_byteenable_2,
	readdata_22,
	readdata_23,
	d_writedata_23,
	readdata_24,
	d_byteenable_3,
	readdata_25,
	readdata_26,
	readdata_4,
	readdata_5,
	d_writedata_14,
	d_byteenable_1,
	readdata_14,
	d_writedata_15,
	readdata_15,
	d_writedata_11,
	readdata_11,
	d_writedata_13,
	readdata_13,
	d_writedata_16,
	readdata_16,
	d_writedata_12,
	readdata_12,
	av_readdata_pre_271,
	av_readdata_pre_281,
	av_readdata_pre_291,
	av_readdata_pre_30,
	av_readdata_pre_311,
	d_writedata_10,
	readdata_10,
	readdata_9,
	readdata_8,
	d_writedata_8,
	readdata_7,
	readdata_6,
	src_payload4,
	d_writedata_21,
	readdata_21,
	d_writedata_20,
	readdata_20,
	src_payload5,
	d_writedata_19,
	readdata_19,
	src_payload6,
	d_writedata_18,
	readdata_18,
	src_payload7,
	d_writedata_17,
	readdata_17,
	src_payload8,
	src_payload9,
	src_payload10,
	src_data_9,
	src_payload11,
	src_payload12,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_32,
	readdata_27,
	readdata_28,
	readdata_29,
	readdata_30,
	readdata_31,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_data_34,
	src_payload24,
	src_payload25,
	src_data_35,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_data_33,
	src_payload31,
	src_payload32,
	src_payload33,
	src_payload34,
	src_payload35,
	src_payload36,
	src_payload37,
	src_payload38,
	src_payload39,
	src_payload40,
	src_payload41,
	src_payload42,
	src_payload43,
	src_payload44,
	src_payload45,
	src_payload46,
	src_payload47,
	src_payload48,
	src_payload49,
	src_payload50,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	sr_0;
output 	W_alu_result_7;
output 	W_alu_result_16;
output 	W_alu_result_15;
output 	W_alu_result_14;
output 	W_alu_result_13;
output 	W_alu_result_12;
output 	W_alu_result_11;
output 	W_alu_result_10;
output 	W_alu_result_9;
output 	W_alu_result_8;
output 	W_alu_result_4;
output 	W_alu_result_5;
output 	W_alu_result_6;
output 	W_alu_result_2;
output 	W_alu_result_3;
input 	q_a_22;
input 	av_readdata_pre_22;
input 	q_a_23;
input 	q_a_24;
input 	q_a_25;
input 	q_a_26;
input 	q_a_1;
input 	q_a_4;
input 	q_a_3;
input 	q_a_2;
input 	q_a_5;
input 	q_a_14;
input 	q_a_15;
input 	q_a_13;
input 	q_a_16;
input 	av_readdata_pre_16;
input 	q_a_12;
input 	q_a_10;
input 	q_a_9;
input 	q_a_8;
input 	q_a_7;
input 	q_a_6;
input 	q_a_21;
input 	av_readdata_pre_21;
input 	q_a_20;
input 	av_readdata_pre_20;
input 	q_a_19;
input 	av_readdata_pre_19;
input 	q_a_18;
input 	av_readdata_pre_18;
input 	q_a_17;
input 	av_readdata_pre_17;
output 	readdata_0;
output 	d_writedata_24;
output 	d_writedata_25;
output 	d_writedata_26;
output 	readdata_1;
output 	readdata_3;
output 	readdata_2;
input 	q_a_27;
input 	q_a_28;
input 	q_a_29;
input 	q_a_30;
input 	q_a_31;
output 	d_writedata_27;
output 	d_writedata_28;
output 	d_writedata_29;
output 	d_writedata_30;
output 	d_writedata_31;
output 	ir_out_0;
output 	ir_out_1;
output 	d_writedata_0;
input 	r_sync_rst;
output 	d_write;
output 	i_read;
output 	F_pc_5;
output 	F_pc_14;
output 	F_pc_13;
output 	F_pc_12;
output 	F_pc_11;
output 	F_pc_10;
output 	F_pc_9;
output 	F_pc_8;
output 	F_pc_7;
output 	F_pc_6;
output 	F_pc_2;
output 	F_pc_3;
output 	F_pc_4;
output 	d_read;
output 	F_pc_1;
output 	F_pc_0;
output 	d_writedata_1;
output 	d_writedata_2;
output 	d_writedata_3;
output 	d_writedata_4;
output 	d_writedata_5;
output 	d_writedata_6;
output 	d_writedata_7;
input 	src0_valid;
input 	read_latency_shift_reg_0;
input 	mem_74_0;
input 	mem_56_0;
input 	src0_valid1;
input 	read_latency_shift_reg_01;
input 	mem_74_01;
input 	mem_56_01;
input 	src0_valid2;
input 	src0_valid3;
input 	WideOr1;
input 	src0_valid4;
input 	read_latency_shift_reg_02;
input 	mem_74_02;
input 	mem_56_02;
input 	src0_valid5;
input 	src0_valid6;
input 	WideOr11;
input 	WideOr12;
input 	saved_grant_0;
output 	debug_mem_slave_waitrequest;
input 	mem_used_1;
input 	av_waitrequest;
input 	src1_valid;
input 	src1_valid1;
input 	src1_valid2;
input 	src1_valid3;
input 	WideOr13;
input 	src1_valid4;
input 	src_payload;
input 	src_payload1;
input 	WideOr14;
input 	uav_write;
output 	d_writedata_9;
input 	WideOr15;
input 	rf_source_valid;
output 	hbreak_enabled;
input 	src_data_0;
input 	av_readdata_pre_221;
input 	av_readdata_pre_23;
input 	av_readdata_pre_24;
input 	av_readdata_pre_25;
input 	av_readdata_pre_26;
input 	src_data_01;
input 	src_data_02;
input 	src_data_03;
input 	av_readdata_pre_1;
input 	av_readdata_pre_11;
input 	av_readdata_pre_12;
input 	av_readdata_pre_13;
input 	av_readdata_pre_14;
input 	av_readdata_pre_15;
input 	av_readdata_pre_4;
input 	av_readdata_pre_41;
input 	av_readdata_pre_42;
input 	av_readdata_pre_43;
input 	av_readdata_pre_3;
input 	src_payload2;
input 	av_readdata_pre_31;
input 	av_readdata_pre_32;
input 	av_readdata_pre_33;
input 	av_readdata_pre_2;
input 	av_readdata_pre_27;
input 	av_readdata_pre_28;
input 	av_readdata_pre_29;
input 	av_readdata_pre_210;
input 	src_data_46;
input 	av_readdata_pre_5;
input 	av_readdata_pre_51;
input 	av_readdata_pre_52;
input 	av_readdata_pre_53;
input 	av_readdata_pre_141;
input 	av_readdata_pre_142;
input 	av_readdata_pre_151;
input 	av_readdata_pre_152;
input 	src_payload3;
input 	av_readdata_pre_111;
input 	av_readdata_pre_131;
input 	av_readdata_pre_132;
input 	av_readdata_pre_161;
input 	av_readdata_pre_121;
input 	av_readdata_pre_122;
input 	av_readdata_pre_10;
input 	av_readdata_pre_101;
input 	av_readdata_pre_9;
input 	av_readdata_pre_91;
input 	av_readdata_pre_92;
input 	av_readdata_pre_8;
input 	av_readdata_pre_81;
input 	av_readdata_pre_82;
input 	av_readdata_pre_7;
input 	av_readdata_pre_71;
input 	av_readdata_pre_72;
input 	av_readdata_pre_73;
input 	av_readdata_pre_6;
input 	av_readdata_pre_61;
input 	av_readdata_pre_62;
input 	av_readdata_pre_63;
input 	av_readdata_pre_211;
input 	av_readdata_pre_201;
input 	av_readdata_pre_191;
input 	av_readdata_pre_181;
input 	av_readdata_pre_171;
input 	r_early_rst;
input 	src_data_8;
output 	d_byteenable_0;
input 	av_readdata_9;
input 	av_readdata_8;
input 	irq;
output 	d_writedata_22;
output 	d_byteenable_2;
output 	readdata_22;
output 	readdata_23;
output 	d_writedata_23;
output 	readdata_24;
output 	d_byteenable_3;
output 	readdata_25;
output 	readdata_26;
output 	readdata_4;
output 	readdata_5;
output 	d_writedata_14;
output 	d_byteenable_1;
output 	readdata_14;
output 	d_writedata_15;
output 	readdata_15;
output 	d_writedata_11;
output 	readdata_11;
output 	d_writedata_13;
output 	readdata_13;
output 	d_writedata_16;
output 	readdata_16;
output 	d_writedata_12;
output 	readdata_12;
input 	av_readdata_pre_271;
input 	av_readdata_pre_281;
input 	av_readdata_pre_291;
input 	av_readdata_pre_30;
input 	av_readdata_pre_311;
output 	d_writedata_10;
output 	readdata_10;
output 	readdata_9;
output 	readdata_8;
output 	d_writedata_8;
output 	readdata_7;
output 	readdata_6;
input 	src_payload4;
output 	d_writedata_21;
output 	readdata_21;
output 	d_writedata_20;
output 	readdata_20;
input 	src_payload5;
output 	d_writedata_19;
output 	readdata_19;
input 	src_payload6;
output 	d_writedata_18;
output 	readdata_18;
input 	src_payload7;
output 	d_writedata_17;
output 	readdata_17;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_data_9;
input 	src_payload11;
input 	src_payload12;
input 	src_data_38;
input 	src_data_39;
input 	src_data_40;
input 	src_data_41;
input 	src_data_42;
input 	src_data_43;
input 	src_data_44;
input 	src_data_45;
input 	src_data_32;
output 	readdata_27;
output 	readdata_28;
output 	readdata_29;
output 	readdata_30;
output 	readdata_31;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_data_34;
input 	src_payload24;
input 	src_payload25;
input 	src_data_35;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_data_33;
input 	src_payload31;
input 	src_payload32;
input 	src_payload33;
input 	src_payload34;
input 	src_payload35;
input 	src_payload36;
input 	src_payload37;
input 	src_payload38;
input 	src_payload39;
input 	src_payload40;
input 	src_payload41;
input 	src_payload42;
input 	src_payload43;
input 	src_payload44;
input 	src_payload45;
input 	src_payload46;
input 	src_payload47;
input 	src_payload48;
input 	src_payload49;
input 	src_payload50;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



processor_processor_nios2_gen2_0_cpu cpu(
	.sr_0(sr_0),
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_16(W_alu_result_16),
	.W_alu_result_15(W_alu_result_15),
	.W_alu_result_14(W_alu_result_14),
	.W_alu_result_13(W_alu_result_13),
	.W_alu_result_12(W_alu_result_12),
	.W_alu_result_11(W_alu_result_11),
	.W_alu_result_10(W_alu_result_10),
	.W_alu_result_9(W_alu_result_9),
	.W_alu_result_8(W_alu_result_8),
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_6(W_alu_result_6),
	.W_alu_result_2(W_alu_result_2),
	.W_alu_result_3(W_alu_result_3),
	.q_a_22(q_a_22),
	.av_readdata_pre_22(av_readdata_pre_22),
	.q_a_23(q_a_23),
	.q_a_24(q_a_24),
	.q_a_25(q_a_25),
	.q_a_26(q_a_26),
	.q_a_1(q_a_1),
	.q_a_4(q_a_4),
	.q_a_3(q_a_3),
	.q_a_2(q_a_2),
	.q_a_5(q_a_5),
	.q_a_14(q_a_14),
	.q_a_15(q_a_15),
	.q_a_13(q_a_13),
	.q_a_16(q_a_16),
	.av_readdata_pre_16(av_readdata_pre_16),
	.q_a_12(q_a_12),
	.q_a_10(q_a_10),
	.q_a_9(q_a_9),
	.q_a_8(q_a_8),
	.q_a_7(q_a_7),
	.q_a_6(q_a_6),
	.q_a_21(q_a_21),
	.av_readdata_pre_21(av_readdata_pre_21),
	.q_a_20(q_a_20),
	.av_readdata_pre_20(av_readdata_pre_20),
	.q_a_19(q_a_19),
	.av_readdata_pre_19(av_readdata_pre_19),
	.q_a_18(q_a_18),
	.av_readdata_pre_18(av_readdata_pre_18),
	.q_a_17(q_a_17),
	.av_readdata_pre_17(av_readdata_pre_17),
	.readdata_0(readdata_0),
	.d_writedata_24(d_writedata_24),
	.d_writedata_25(d_writedata_25),
	.d_writedata_26(d_writedata_26),
	.readdata_1(readdata_1),
	.readdata_3(readdata_3),
	.readdata_2(readdata_2),
	.q_a_27(q_a_27),
	.q_a_28(q_a_28),
	.q_a_29(q_a_29),
	.q_a_30(q_a_30),
	.q_a_31(q_a_31),
	.d_writedata_27(d_writedata_27),
	.d_writedata_28(d_writedata_28),
	.d_writedata_29(d_writedata_29),
	.d_writedata_30(d_writedata_30),
	.d_writedata_31(d_writedata_31),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.d_writedata_0(d_writedata_0),
	.r_sync_rst(r_sync_rst),
	.d_write1(d_write),
	.i_read1(i_read),
	.F_pc_5(F_pc_5),
	.F_pc_14(F_pc_14),
	.F_pc_13(F_pc_13),
	.F_pc_12(F_pc_12),
	.F_pc_11(F_pc_11),
	.F_pc_10(F_pc_10),
	.F_pc_9(F_pc_9),
	.F_pc_8(F_pc_8),
	.F_pc_7(F_pc_7),
	.F_pc_6(F_pc_6),
	.F_pc_2(F_pc_2),
	.F_pc_3(F_pc_3),
	.F_pc_4(F_pc_4),
	.d_read1(d_read),
	.F_pc_1(F_pc_1),
	.F_pc_0(F_pc_0),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.src0_valid(src0_valid),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.mem_74_0(mem_74_0),
	.mem_56_0(mem_56_0),
	.src0_valid1(src0_valid1),
	.read_latency_shift_reg_01(read_latency_shift_reg_01),
	.mem_74_01(mem_74_01),
	.mem_56_01(mem_56_01),
	.src0_valid2(src0_valid2),
	.src0_valid3(src0_valid3),
	.WideOr1(WideOr1),
	.src0_valid4(src0_valid4),
	.read_latency_shift_reg_02(read_latency_shift_reg_02),
	.mem_74_02(mem_74_02),
	.mem_56_02(mem_56_02),
	.src0_valid5(src0_valid5),
	.src0_valid6(src0_valid6),
	.WideOr11(WideOr11),
	.WideOr12(WideOr12),
	.saved_grant_0(saved_grant_0),
	.debug_mem_slave_waitrequest(debug_mem_slave_waitrequest),
	.mem_used_1(mem_used_1),
	.av_waitrequest(av_waitrequest),
	.src1_valid(src1_valid),
	.src1_valid1(src1_valid1),
	.src1_valid2(src1_valid2),
	.src1_valid3(src1_valid3),
	.WideOr13(WideOr13),
	.src1_valid4(src1_valid4),
	.src_payload(src_payload),
	.src_payload1(src_payload1),
	.WideOr14(WideOr14),
	.uav_write(uav_write),
	.d_writedata_9(d_writedata_9),
	.WideOr15(WideOr15),
	.rf_source_valid(rf_source_valid),
	.hbreak_enabled1(hbreak_enabled),
	.src_data_0(src_data_0),
	.av_readdata_pre_221(av_readdata_pre_221),
	.av_readdata_pre_23(av_readdata_pre_23),
	.av_readdata_pre_24(av_readdata_pre_24),
	.av_readdata_pre_25(av_readdata_pre_25),
	.av_readdata_pre_26(av_readdata_pre_26),
	.src_data_01(src_data_01),
	.src_data_02(src_data_02),
	.src_data_03(src_data_03),
	.av_readdata_pre_1(av_readdata_pre_1),
	.av_readdata_pre_11(av_readdata_pre_11),
	.av_readdata_pre_12(av_readdata_pre_12),
	.av_readdata_pre_13(av_readdata_pre_13),
	.av_readdata_pre_14(av_readdata_pre_14),
	.av_readdata_pre_15(av_readdata_pre_15),
	.av_readdata_pre_4(av_readdata_pre_4),
	.av_readdata_pre_41(av_readdata_pre_41),
	.av_readdata_pre_42(av_readdata_pre_42),
	.av_readdata_pre_43(av_readdata_pre_43),
	.av_readdata_pre_3(av_readdata_pre_3),
	.src_payload2(src_payload2),
	.av_readdata_pre_31(av_readdata_pre_31),
	.av_readdata_pre_32(av_readdata_pre_32),
	.av_readdata_pre_33(av_readdata_pre_33),
	.av_readdata_pre_2(av_readdata_pre_2),
	.av_readdata_pre_27(av_readdata_pre_27),
	.av_readdata_pre_28(av_readdata_pre_28),
	.av_readdata_pre_29(av_readdata_pre_29),
	.av_readdata_pre_210(av_readdata_pre_210),
	.src_data_46(src_data_46),
	.av_readdata_pre_5(av_readdata_pre_5),
	.av_readdata_pre_51(av_readdata_pre_51),
	.av_readdata_pre_52(av_readdata_pre_52),
	.av_readdata_pre_53(av_readdata_pre_53),
	.av_readdata_pre_141(av_readdata_pre_141),
	.av_readdata_pre_142(av_readdata_pre_142),
	.av_readdata_pre_151(av_readdata_pre_151),
	.av_readdata_pre_152(av_readdata_pre_152),
	.src_payload3(src_payload3),
	.av_readdata_pre_111(av_readdata_pre_111),
	.av_readdata_pre_131(av_readdata_pre_131),
	.av_readdata_pre_132(av_readdata_pre_132),
	.av_readdata_pre_161(av_readdata_pre_161),
	.av_readdata_pre_121(av_readdata_pre_121),
	.av_readdata_pre_122(av_readdata_pre_122),
	.av_readdata_pre_10(av_readdata_pre_10),
	.av_readdata_pre_101(av_readdata_pre_101),
	.av_readdata_pre_9(av_readdata_pre_9),
	.av_readdata_pre_91(av_readdata_pre_91),
	.av_readdata_pre_92(av_readdata_pre_92),
	.av_readdata_pre_8(av_readdata_pre_8),
	.av_readdata_pre_81(av_readdata_pre_81),
	.av_readdata_pre_82(av_readdata_pre_82),
	.av_readdata_pre_7(av_readdata_pre_7),
	.av_readdata_pre_71(av_readdata_pre_71),
	.av_readdata_pre_72(av_readdata_pre_72),
	.av_readdata_pre_73(av_readdata_pre_73),
	.av_readdata_pre_6(av_readdata_pre_6),
	.av_readdata_pre_61(av_readdata_pre_61),
	.av_readdata_pre_62(av_readdata_pre_62),
	.av_readdata_pre_63(av_readdata_pre_63),
	.av_readdata_pre_211(av_readdata_pre_211),
	.av_readdata_pre_201(av_readdata_pre_201),
	.av_readdata_pre_191(av_readdata_pre_191),
	.av_readdata_pre_181(av_readdata_pre_181),
	.av_readdata_pre_171(av_readdata_pre_171),
	.r_early_rst(r_early_rst),
	.src_data_8(src_data_8),
	.d_byteenable_0(d_byteenable_0),
	.av_readdata_9(av_readdata_9),
	.av_readdata_8(av_readdata_8),
	.irq(irq),
	.d_writedata_22(d_writedata_22),
	.d_byteenable_2(d_byteenable_2),
	.readdata_22(readdata_22),
	.readdata_23(readdata_23),
	.d_writedata_23(d_writedata_23),
	.readdata_24(readdata_24),
	.d_byteenable_3(d_byteenable_3),
	.readdata_25(readdata_25),
	.readdata_26(readdata_26),
	.readdata_4(readdata_4),
	.readdata_5(readdata_5),
	.d_writedata_14(d_writedata_14),
	.d_byteenable_1(d_byteenable_1),
	.readdata_14(readdata_14),
	.d_writedata_15(d_writedata_15),
	.readdata_15(readdata_15),
	.d_writedata_11(d_writedata_11),
	.readdata_11(readdata_11),
	.d_writedata_13(d_writedata_13),
	.readdata_13(readdata_13),
	.d_writedata_16(d_writedata_16),
	.readdata_16(readdata_16),
	.d_writedata_12(d_writedata_12),
	.readdata_12(readdata_12),
	.av_readdata_pre_271(av_readdata_pre_271),
	.av_readdata_pre_281(av_readdata_pre_281),
	.av_readdata_pre_291(av_readdata_pre_291),
	.av_readdata_pre_30(av_readdata_pre_30),
	.av_readdata_pre_311(av_readdata_pre_311),
	.d_writedata_10(d_writedata_10),
	.readdata_10(readdata_10),
	.readdata_9(readdata_9),
	.readdata_8(readdata_8),
	.d_writedata_8(d_writedata_8),
	.readdata_7(readdata_7),
	.readdata_6(readdata_6),
	.src_payload4(src_payload4),
	.d_writedata_21(d_writedata_21),
	.readdata_21(readdata_21),
	.d_writedata_20(d_writedata_20),
	.readdata_20(readdata_20),
	.src_payload5(src_payload5),
	.d_writedata_19(d_writedata_19),
	.readdata_19(readdata_19),
	.src_payload6(src_payload6),
	.d_writedata_18(d_writedata_18),
	.readdata_18(readdata_18),
	.src_payload7(src_payload7),
	.d_writedata_17(d_writedata_17),
	.readdata_17(readdata_17),
	.src_payload8(src_payload8),
	.src_payload9(src_payload9),
	.src_payload10(src_payload10),
	.src_data_9(src_data_9),
	.src_payload11(src_payload11),
	.src_payload12(src_payload12),
	.src_data_38(src_data_38),
	.src_data_39(src_data_39),
	.src_data_40(src_data_40),
	.src_data_41(src_data_41),
	.src_data_42(src_data_42),
	.src_data_43(src_data_43),
	.src_data_44(src_data_44),
	.src_data_45(src_data_45),
	.src_data_32(src_data_32),
	.readdata_27(readdata_27),
	.readdata_28(readdata_28),
	.readdata_29(readdata_29),
	.readdata_30(readdata_30),
	.readdata_31(readdata_31),
	.src_payload13(src_payload13),
	.src_payload14(src_payload14),
	.src_payload15(src_payload15),
	.src_payload16(src_payload16),
	.src_payload17(src_payload17),
	.src_payload18(src_payload18),
	.src_payload19(src_payload19),
	.src_payload20(src_payload20),
	.src_payload21(src_payload21),
	.src_payload22(src_payload22),
	.src_payload23(src_payload23),
	.src_data_34(src_data_34),
	.src_payload24(src_payload24),
	.src_payload25(src_payload25),
	.src_data_35(src_data_35),
	.src_payload26(src_payload26),
	.src_payload27(src_payload27),
	.src_payload28(src_payload28),
	.src_payload29(src_payload29),
	.src_payload30(src_payload30),
	.src_data_33(src_data_33),
	.src_payload31(src_payload31),
	.src_payload32(src_payload32),
	.src_payload33(src_payload33),
	.src_payload34(src_payload34),
	.src_payload35(src_payload35),
	.src_payload36(src_payload36),
	.src_payload37(src_payload37),
	.src_payload38(src_payload38),
	.src_payload39(src_payload39),
	.src_payload40(src_payload40),
	.src_payload41(src_payload41),
	.src_payload42(src_payload42),
	.src_payload43(src_payload43),
	.src_payload44(src_payload44),
	.src_payload45(src_payload45),
	.src_payload46(src_payload46),
	.src_payload47(src_payload47),
	.src_payload48(src_payload48),
	.src_payload49(src_payload49),
	.src_payload50(src_payload50),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_1(state_1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2),
	.clk_clk(clk_clk));

endmodule

module processor_processor_nios2_gen2_0_cpu (
	sr_0,
	W_alu_result_7,
	W_alu_result_16,
	W_alu_result_15,
	W_alu_result_14,
	W_alu_result_13,
	W_alu_result_12,
	W_alu_result_11,
	W_alu_result_10,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_4,
	W_alu_result_5,
	W_alu_result_6,
	W_alu_result_2,
	W_alu_result_3,
	q_a_22,
	av_readdata_pre_22,
	q_a_23,
	q_a_24,
	q_a_25,
	q_a_26,
	q_a_1,
	q_a_4,
	q_a_3,
	q_a_2,
	q_a_5,
	q_a_14,
	q_a_15,
	q_a_13,
	q_a_16,
	av_readdata_pre_16,
	q_a_12,
	q_a_10,
	q_a_9,
	q_a_8,
	q_a_7,
	q_a_6,
	q_a_21,
	av_readdata_pre_21,
	q_a_20,
	av_readdata_pre_20,
	q_a_19,
	av_readdata_pre_19,
	q_a_18,
	av_readdata_pre_18,
	q_a_17,
	av_readdata_pre_17,
	readdata_0,
	d_writedata_24,
	d_writedata_25,
	d_writedata_26,
	readdata_1,
	readdata_3,
	readdata_2,
	q_a_27,
	q_a_28,
	q_a_29,
	q_a_30,
	q_a_31,
	d_writedata_27,
	d_writedata_28,
	d_writedata_29,
	d_writedata_30,
	d_writedata_31,
	ir_out_0,
	ir_out_1,
	d_writedata_0,
	r_sync_rst,
	d_write1,
	i_read1,
	F_pc_5,
	F_pc_14,
	F_pc_13,
	F_pc_12,
	F_pc_11,
	F_pc_10,
	F_pc_9,
	F_pc_8,
	F_pc_7,
	F_pc_6,
	F_pc_2,
	F_pc_3,
	F_pc_4,
	d_read1,
	F_pc_1,
	F_pc_0,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	src0_valid,
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	src0_valid1,
	read_latency_shift_reg_01,
	mem_74_01,
	mem_56_01,
	src0_valid2,
	src0_valid3,
	WideOr1,
	src0_valid4,
	read_latency_shift_reg_02,
	mem_74_02,
	mem_56_02,
	src0_valid5,
	src0_valid6,
	WideOr11,
	WideOr12,
	saved_grant_0,
	debug_mem_slave_waitrequest,
	mem_used_1,
	av_waitrequest,
	src1_valid,
	src1_valid1,
	src1_valid2,
	src1_valid3,
	WideOr13,
	src1_valid4,
	src_payload,
	src_payload1,
	WideOr14,
	uav_write,
	d_writedata_9,
	WideOr15,
	rf_source_valid,
	hbreak_enabled1,
	src_data_0,
	av_readdata_pre_221,
	av_readdata_pre_23,
	av_readdata_pre_24,
	av_readdata_pre_25,
	av_readdata_pre_26,
	src_data_01,
	src_data_02,
	src_data_03,
	av_readdata_pre_1,
	av_readdata_pre_11,
	av_readdata_pre_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	av_readdata_pre_15,
	av_readdata_pre_4,
	av_readdata_pre_41,
	av_readdata_pre_42,
	av_readdata_pre_43,
	av_readdata_pre_3,
	src_payload2,
	av_readdata_pre_31,
	av_readdata_pre_32,
	av_readdata_pre_33,
	av_readdata_pre_2,
	av_readdata_pre_27,
	av_readdata_pre_28,
	av_readdata_pre_29,
	av_readdata_pre_210,
	src_data_46,
	av_readdata_pre_5,
	av_readdata_pre_51,
	av_readdata_pre_52,
	av_readdata_pre_53,
	av_readdata_pre_141,
	av_readdata_pre_142,
	av_readdata_pre_151,
	av_readdata_pre_152,
	src_payload3,
	av_readdata_pre_111,
	av_readdata_pre_131,
	av_readdata_pre_132,
	av_readdata_pre_161,
	av_readdata_pre_121,
	av_readdata_pre_122,
	av_readdata_pre_10,
	av_readdata_pre_101,
	av_readdata_pre_9,
	av_readdata_pre_91,
	av_readdata_pre_92,
	av_readdata_pre_8,
	av_readdata_pre_81,
	av_readdata_pre_82,
	av_readdata_pre_7,
	av_readdata_pre_71,
	av_readdata_pre_72,
	av_readdata_pre_73,
	av_readdata_pre_6,
	av_readdata_pre_61,
	av_readdata_pre_62,
	av_readdata_pre_63,
	av_readdata_pre_211,
	av_readdata_pre_201,
	av_readdata_pre_191,
	av_readdata_pre_181,
	av_readdata_pre_171,
	r_early_rst,
	src_data_8,
	d_byteenable_0,
	av_readdata_9,
	av_readdata_8,
	irq,
	d_writedata_22,
	d_byteenable_2,
	readdata_22,
	readdata_23,
	d_writedata_23,
	readdata_24,
	d_byteenable_3,
	readdata_25,
	readdata_26,
	readdata_4,
	readdata_5,
	d_writedata_14,
	d_byteenable_1,
	readdata_14,
	d_writedata_15,
	readdata_15,
	d_writedata_11,
	readdata_11,
	d_writedata_13,
	readdata_13,
	d_writedata_16,
	readdata_16,
	d_writedata_12,
	readdata_12,
	av_readdata_pre_271,
	av_readdata_pre_281,
	av_readdata_pre_291,
	av_readdata_pre_30,
	av_readdata_pre_311,
	d_writedata_10,
	readdata_10,
	readdata_9,
	readdata_8,
	d_writedata_8,
	readdata_7,
	readdata_6,
	src_payload4,
	d_writedata_21,
	readdata_21,
	d_writedata_20,
	readdata_20,
	src_payload5,
	d_writedata_19,
	readdata_19,
	src_payload6,
	d_writedata_18,
	readdata_18,
	src_payload7,
	d_writedata_17,
	readdata_17,
	src_payload8,
	src_payload9,
	src_payload10,
	src_data_9,
	src_payload11,
	src_payload12,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_32,
	readdata_27,
	readdata_28,
	readdata_29,
	readdata_30,
	readdata_31,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_data_34,
	src_payload24,
	src_payload25,
	src_data_35,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_data_33,
	src_payload31,
	src_payload32,
	src_payload33,
	src_payload34,
	src_payload35,
	src_payload36,
	src_payload37,
	src_payload38,
	src_payload39,
	src_payload40,
	src_payload41,
	src_payload42,
	src_payload43,
	src_payload44,
	src_payload45,
	src_payload46,
	src_payload47,
	src_payload48,
	src_payload49,
	src_payload50,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	sr_0;
output 	W_alu_result_7;
output 	W_alu_result_16;
output 	W_alu_result_15;
output 	W_alu_result_14;
output 	W_alu_result_13;
output 	W_alu_result_12;
output 	W_alu_result_11;
output 	W_alu_result_10;
output 	W_alu_result_9;
output 	W_alu_result_8;
output 	W_alu_result_4;
output 	W_alu_result_5;
output 	W_alu_result_6;
output 	W_alu_result_2;
output 	W_alu_result_3;
input 	q_a_22;
input 	av_readdata_pre_22;
input 	q_a_23;
input 	q_a_24;
input 	q_a_25;
input 	q_a_26;
input 	q_a_1;
input 	q_a_4;
input 	q_a_3;
input 	q_a_2;
input 	q_a_5;
input 	q_a_14;
input 	q_a_15;
input 	q_a_13;
input 	q_a_16;
input 	av_readdata_pre_16;
input 	q_a_12;
input 	q_a_10;
input 	q_a_9;
input 	q_a_8;
input 	q_a_7;
input 	q_a_6;
input 	q_a_21;
input 	av_readdata_pre_21;
input 	q_a_20;
input 	av_readdata_pre_20;
input 	q_a_19;
input 	av_readdata_pre_19;
input 	q_a_18;
input 	av_readdata_pre_18;
input 	q_a_17;
input 	av_readdata_pre_17;
output 	readdata_0;
output 	d_writedata_24;
output 	d_writedata_25;
output 	d_writedata_26;
output 	readdata_1;
output 	readdata_3;
output 	readdata_2;
input 	q_a_27;
input 	q_a_28;
input 	q_a_29;
input 	q_a_30;
input 	q_a_31;
output 	d_writedata_27;
output 	d_writedata_28;
output 	d_writedata_29;
output 	d_writedata_30;
output 	d_writedata_31;
output 	ir_out_0;
output 	ir_out_1;
output 	d_writedata_0;
input 	r_sync_rst;
output 	d_write1;
output 	i_read1;
output 	F_pc_5;
output 	F_pc_14;
output 	F_pc_13;
output 	F_pc_12;
output 	F_pc_11;
output 	F_pc_10;
output 	F_pc_9;
output 	F_pc_8;
output 	F_pc_7;
output 	F_pc_6;
output 	F_pc_2;
output 	F_pc_3;
output 	F_pc_4;
output 	d_read1;
output 	F_pc_1;
output 	F_pc_0;
output 	d_writedata_1;
output 	d_writedata_2;
output 	d_writedata_3;
output 	d_writedata_4;
output 	d_writedata_5;
output 	d_writedata_6;
output 	d_writedata_7;
input 	src0_valid;
input 	read_latency_shift_reg_0;
input 	mem_74_0;
input 	mem_56_0;
input 	src0_valid1;
input 	read_latency_shift_reg_01;
input 	mem_74_01;
input 	mem_56_01;
input 	src0_valid2;
input 	src0_valid3;
input 	WideOr1;
input 	src0_valid4;
input 	read_latency_shift_reg_02;
input 	mem_74_02;
input 	mem_56_02;
input 	src0_valid5;
input 	src0_valid6;
input 	WideOr11;
input 	WideOr12;
input 	saved_grant_0;
output 	debug_mem_slave_waitrequest;
input 	mem_used_1;
input 	av_waitrequest;
input 	src1_valid;
input 	src1_valid1;
input 	src1_valid2;
input 	src1_valid3;
input 	WideOr13;
input 	src1_valid4;
input 	src_payload;
input 	src_payload1;
input 	WideOr14;
input 	uav_write;
output 	d_writedata_9;
input 	WideOr15;
input 	rf_source_valid;
output 	hbreak_enabled1;
input 	src_data_0;
input 	av_readdata_pre_221;
input 	av_readdata_pre_23;
input 	av_readdata_pre_24;
input 	av_readdata_pre_25;
input 	av_readdata_pre_26;
input 	src_data_01;
input 	src_data_02;
input 	src_data_03;
input 	av_readdata_pre_1;
input 	av_readdata_pre_11;
input 	av_readdata_pre_12;
input 	av_readdata_pre_13;
input 	av_readdata_pre_14;
input 	av_readdata_pre_15;
input 	av_readdata_pre_4;
input 	av_readdata_pre_41;
input 	av_readdata_pre_42;
input 	av_readdata_pre_43;
input 	av_readdata_pre_3;
input 	src_payload2;
input 	av_readdata_pre_31;
input 	av_readdata_pre_32;
input 	av_readdata_pre_33;
input 	av_readdata_pre_2;
input 	av_readdata_pre_27;
input 	av_readdata_pre_28;
input 	av_readdata_pre_29;
input 	av_readdata_pre_210;
input 	src_data_46;
input 	av_readdata_pre_5;
input 	av_readdata_pre_51;
input 	av_readdata_pre_52;
input 	av_readdata_pre_53;
input 	av_readdata_pre_141;
input 	av_readdata_pre_142;
input 	av_readdata_pre_151;
input 	av_readdata_pre_152;
input 	src_payload3;
input 	av_readdata_pre_111;
input 	av_readdata_pre_131;
input 	av_readdata_pre_132;
input 	av_readdata_pre_161;
input 	av_readdata_pre_121;
input 	av_readdata_pre_122;
input 	av_readdata_pre_10;
input 	av_readdata_pre_101;
input 	av_readdata_pre_9;
input 	av_readdata_pre_91;
input 	av_readdata_pre_92;
input 	av_readdata_pre_8;
input 	av_readdata_pre_81;
input 	av_readdata_pre_82;
input 	av_readdata_pre_7;
input 	av_readdata_pre_71;
input 	av_readdata_pre_72;
input 	av_readdata_pre_73;
input 	av_readdata_pre_6;
input 	av_readdata_pre_61;
input 	av_readdata_pre_62;
input 	av_readdata_pre_63;
input 	av_readdata_pre_211;
input 	av_readdata_pre_201;
input 	av_readdata_pre_191;
input 	av_readdata_pre_181;
input 	av_readdata_pre_171;
input 	r_early_rst;
input 	src_data_8;
output 	d_byteenable_0;
input 	av_readdata_9;
input 	av_readdata_8;
input 	irq;
output 	d_writedata_22;
output 	d_byteenable_2;
output 	readdata_22;
output 	readdata_23;
output 	d_writedata_23;
output 	readdata_24;
output 	d_byteenable_3;
output 	readdata_25;
output 	readdata_26;
output 	readdata_4;
output 	readdata_5;
output 	d_writedata_14;
output 	d_byteenable_1;
output 	readdata_14;
output 	d_writedata_15;
output 	readdata_15;
output 	d_writedata_11;
output 	readdata_11;
output 	d_writedata_13;
output 	readdata_13;
output 	d_writedata_16;
output 	readdata_16;
output 	d_writedata_12;
output 	readdata_12;
input 	av_readdata_pre_271;
input 	av_readdata_pre_281;
input 	av_readdata_pre_291;
input 	av_readdata_pre_30;
input 	av_readdata_pre_311;
output 	d_writedata_10;
output 	readdata_10;
output 	readdata_9;
output 	readdata_8;
output 	d_writedata_8;
output 	readdata_7;
output 	readdata_6;
input 	src_payload4;
output 	d_writedata_21;
output 	readdata_21;
output 	d_writedata_20;
output 	readdata_20;
input 	src_payload5;
output 	d_writedata_19;
output 	readdata_19;
input 	src_payload6;
output 	d_writedata_18;
output 	readdata_18;
input 	src_payload7;
output 	d_writedata_17;
output 	readdata_17;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_data_9;
input 	src_payload11;
input 	src_payload12;
input 	src_data_38;
input 	src_data_39;
input 	src_data_40;
input 	src_data_41;
input 	src_data_42;
input 	src_data_43;
input 	src_data_44;
input 	src_data_45;
input 	src_data_32;
output 	readdata_27;
output 	readdata_28;
output 	readdata_29;
output 	readdata_30;
output 	readdata_31;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_data_34;
input 	src_payload24;
input 	src_payload25;
input 	src_data_35;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_data_33;
input 	src_payload31;
input 	src_payload32;
input 	src_payload33;
input 	src_payload34;
input 	src_payload35;
input 	src_payload36;
input 	src_payload37;
input 	src_payload38;
input 	src_payload39;
input 	src_payload40;
input 	src_payload41;
input 	src_payload42;
input 	src_payload43;
input 	src_payload44;
input 	src_payload45;
input 	src_payload46;
input 	src_payload47;
input 	src_payload48;
input 	src_payload49;
input 	src_payload50;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ;
wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ;
wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ;
wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ;
wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ;
wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ;
wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ;
wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ;
wire \W_alu_result[0]~q ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[7] ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[6] ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[5] ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[4] ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[3] ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[2] ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[1] ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[0] ;
wire \Add1~68_combout ;
wire \Add1~70_combout ;
wire \Add1~72_combout ;
wire \Add1~74_combout ;
wire \Add1~76_combout ;
wire \Add1~78_combout ;
wire \Add1~80_combout ;
wire \Add1~82_combout ;
wire \Add1~84_combout ;
wire \Add1~86_combout ;
wire \Add1~88_combout ;
wire \Add1~90_combout ;
wire \Add1~92_combout ;
wire \Add1~94_combout ;
wire \Add1~96_combout ;
wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[16] ;
wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[15] ;
wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[14] ;
wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[13] ;
wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[12] ;
wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[11] ;
wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[10] ;
wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[9] ;
wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[8] ;
wire \W_alu_result[1]~q ;
wire \av_ld_byte1_data[0]~q ;
wire \W_alu_result[0]~15_combout ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci|the_processor_nios2_gen2_0_cpu_nios2_oci_debug|jtag_break~q ;
wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[31] ;
wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[30] ;
wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[29] ;
wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[28] ;
wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[27] ;
wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[26] ;
wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[25] ;
wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[24] ;
wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[23] ;
wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[22] ;
wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[21] ;
wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[20] ;
wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[19] ;
wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[18] ;
wire \processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ;
wire \processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[17] ;
wire \av_ld_byte2_data[0]~q ;
wire \av_ld_byte1_data[7]~q ;
wire \av_ld_byte1_data[6]~q ;
wire \av_ld_byte1_data[5]~q ;
wire \av_ld_byte1_data[4]~q ;
wire \av_ld_byte1_data[3]~q ;
wire \av_ld_byte1_data[2]~q ;
wire \av_ld_byte1_data[1]~q ;
wire \W_alu_result[1]~16_combout ;
wire \av_ld_byte1_data[0]~0_combout ;
wire \W_alu_result[31]~q ;
wire \W_alu_result[30]~q ;
wire \W_alu_result[29]~q ;
wire \W_alu_result[28]~q ;
wire \W_alu_result[27]~q ;
wire \W_alu_result[26]~q ;
wire \W_alu_result[25]~q ;
wire \W_alu_result[24]~q ;
wire \av_ld_byte2_data[7]~q ;
wire \W_alu_result[23]~q ;
wire \av_ld_byte2_data[6]~q ;
wire \W_alu_result[22]~q ;
wire \av_ld_byte2_data[5]~q ;
wire \W_alu_result[21]~q ;
wire \av_ld_byte2_data[4]~q ;
wire \W_alu_result[20]~q ;
wire \av_ld_byte2_data[3]~q ;
wire \W_alu_result[19]~q ;
wire \av_ld_byte2_data[2]~q ;
wire \W_alu_result[18]~q ;
wire \av_ld_byte2_data[1]~q ;
wire \W_alu_result[17]~q ;
wire \av_ld_byte2_data[0]~0_combout ;
wire \av_ld_byte1_data[7]~1_combout ;
wire \av_ld_byte1_data[6]~2_combout ;
wire \av_ld_byte1_data[5]~3_combout ;
wire \av_ld_byte1_data[4]~4_combout ;
wire \av_ld_byte1_data[3]~5_combout ;
wire \av_ld_byte1_data[2]~6_combout ;
wire \av_ld_byte1_data[1]~7_combout ;
wire \W_alu_result[31]~17_combout ;
wire \W_alu_result[30]~18_combout ;
wire \W_alu_result[29]~31_combout ;
wire \W_alu_result[28]~19_combout ;
wire \W_alu_result[27]~20_combout ;
wire \W_alu_result[26]~21_combout ;
wire \W_alu_result[25]~22_combout ;
wire \W_alu_result[24]~23_combout ;
wire \av_ld_byte2_data[7]~1_combout ;
wire \W_alu_result[23]~24_combout ;
wire \av_ld_byte2_data[6]~2_combout ;
wire \W_alu_result[22]~25_combout ;
wire \av_ld_byte2_data[5]~3_combout ;
wire \W_alu_result[21]~26_combout ;
wire \av_ld_byte2_data[4]~4_combout ;
wire \W_alu_result[20]~27_combout ;
wire \av_ld_byte2_data[3]~5_combout ;
wire \W_alu_result[19]~28_combout ;
wire \av_ld_byte2_data[2]~6_combout ;
wire \W_alu_result[18]~29_combout ;
wire \av_ld_byte2_data[1]~7_combout ;
wire \W_alu_result[17]~30_combout ;
wire \R_wr_dst_reg~q ;
wire \W_rf_wren~combout ;
wire \av_ld_byte0_data[0]~q ;
wire \W_rf_wr_data[0]~0_combout ;
wire \W_control_rd_data[0]~q ;
wire \W_rf_wr_data[0]~1_combout ;
wire \W_rf_wr_data[0]~2_combout ;
wire \R_dst_regnum[0]~q ;
wire \R_dst_regnum[1]~q ;
wire \R_dst_regnum[2]~q ;
wire \R_dst_regnum[3]~q ;
wire \R_dst_regnum[4]~q ;
wire \D_iw[22]~q ;
wire \D_iw[23]~q ;
wire \D_iw[24]~q ;
wire \D_iw[25]~q ;
wire \D_iw[26]~q ;
wire \D_ctrl_ld_signed~1_combout ;
wire \av_ld_byte0_data[1]~q ;
wire \W_control_rd_data[1]~q ;
wire \W_rf_wr_data[1]~3_combout ;
wire \W_rf_wr_data[1]~4_combout ;
wire \av_ld_byte0_data[2]~q ;
wire \W_rf_wr_data[2]~5_combout ;
wire \av_ld_byte0_data[3]~q ;
wire \W_rf_wr_data[3]~6_combout ;
wire \av_ld_byte0_data[4]~q ;
wire \W_rf_wr_data[4]~7_combout ;
wire \av_ld_byte0_data[5]~q ;
wire \W_rf_wr_data[5]~8_combout ;
wire \av_ld_byte0_data[6]~q ;
wire \W_rf_wr_data[6]~9_combout ;
wire \av_ld_byte0_data[7]~q ;
wire \W_rf_wr_data[7]~10_combout ;
wire \D_wr_dst_reg~0_combout ;
wire \D_wr_dst_reg~1_combout ;
wire \D_ctrl_implicit_dst_eretaddr~5_combout ;
wire \D_ctrl_implicit_dst_eretaddr~6_combout ;
wire \D_ctrl_implicit_dst_eretaddr~7_combout ;
wire \D_ctrl_implicit_dst_eretaddr~8_combout ;
wire \D_dst_regnum[0]~2_combout ;
wire \D_dst_regnum[1]~3_combout ;
wire \D_dst_regnum[0]~4_combout ;
wire \Equal0~19_combout ;
wire \D_dst_regnum[3]~5_combout ;
wire \D_dst_regnum[4]~6_combout ;
wire \Equal0~20_combout ;
wire \D_dst_regnum[2]~7_combout ;
wire \D_wr_dst_reg~2_combout ;
wire \av_ld_rshift8~0_combout ;
wire \av_ld_rshift8~1_combout ;
wire \av_ld_byte0_data[7]~0_combout ;
wire \E_control_rd_data[0]~0_combout ;
wire \E_control_rd_data[0]~1_combout ;
wire \E_control_rd_data[0]~2_combout ;
wire \E_control_rd_data[0]~3_combout ;
wire \D_dst_regnum[0]~8_combout ;
wire \D_dst_regnum[3]~9_combout ;
wire \D_dst_regnum[4]~10_combout ;
wire \F_iw[22]~4_combout ;
wire \F_iw[22]~5_combout ;
wire \F_iw[23]~6_combout ;
wire \F_iw[23]~7_combout ;
wire \F_iw[24]~8_combout ;
wire \F_iw[24]~9_combout ;
wire \F_iw[25]~10_combout ;
wire \F_iw[25]~11_combout ;
wire \F_iw[26]~12_combout ;
wire \F_iw[26]~13_combout ;
wire \D_iw[27]~q ;
wire \D_iw[28]~q ;
wire \D_iw[29]~q ;
wire \D_iw[30]~q ;
wire \D_iw[31]~q ;
wire \W_rf_wr_data[16]~11_combout ;
wire \W_rf_wr_data[15]~12_combout ;
wire \W_rf_wr_data[14]~13_combout ;
wire \W_rf_wr_data[13]~14_combout ;
wire \W_rf_wr_data[12]~15_combout ;
wire \W_rf_wr_data[11]~16_combout ;
wire \W_rf_wr_data[10]~17_combout ;
wire \W_rf_wr_data[9]~18_combout ;
wire \W_rf_wr_data[8]~19_combout ;
wire \av_ld_byte0_data_nxt[1]~12_combout ;
wire \av_ld_byte0_data_nxt[1]~13_combout ;
wire \av_ld_byte0_data_nxt[1]~14_combout ;
wire \av_ld_byte0_data_nxt[1]~15_combout ;
wire \av_ld_byte0_data_nxt[1]~16_combout ;
wire \av_ld_byte0_data_nxt[1]~17_combout ;
wire \E_control_rd_data[1]~4_combout ;
wire \E_control_rd_data[1]~5_combout ;
wire \av_ld_byte0_data_nxt[2]~18_combout ;
wire \av_ld_byte0_data_nxt[2]~19_combout ;
wire \av_ld_byte0_data_nxt[2]~20_combout ;
wire \av_ld_byte0_data_nxt[2]~21_combout ;
wire \av_ld_byte0_data_nxt[2]~22_combout ;
wire \av_ld_byte0_data_nxt[3]~23_combout ;
wire \av_ld_byte0_data_nxt[3]~24_combout ;
wire \av_ld_byte0_data_nxt[3]~25_combout ;
wire \av_ld_byte0_data_nxt[4]~26_combout ;
wire \av_ld_byte0_data_nxt[4]~27_combout ;
wire \av_ld_byte0_data_nxt[4]~28_combout ;
wire \av_ld_byte0_data_nxt[5]~29_combout ;
wire \av_ld_byte0_data_nxt[5]~30_combout ;
wire \av_ld_byte0_data_nxt[5]~31_combout ;
wire \av_ld_byte0_data_nxt[6]~32_combout ;
wire \av_ld_byte0_data_nxt[6]~33_combout ;
wire \av_ld_byte0_data_nxt[6]~34_combout ;
wire \av_ld_byte0_data_nxt[7]~35_combout ;
wire \av_ld_byte0_data_nxt[7]~36_combout ;
wire \av_ld_byte0_data_nxt[7]~37_combout ;
wire \R_ctrl_ld_signed~q ;
wire \av_fill_bit~0_combout ;
wire \av_ld_byte1_data_en~0_combout ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci|the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[0]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci|the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[1]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci|the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_single_step_mode~q ;
wire \F_iw[27]~73_combout ;
wire \F_iw[27]~74_combout ;
wire \F_iw[28]~75_combout ;
wire \F_iw[28]~76_combout ;
wire \F_iw[29]~77_combout ;
wire \F_iw[29]~78_combout ;
wire \F_iw[30]~79_combout ;
wire \F_iw[30]~80_combout ;
wire \F_iw[31]~81_combout ;
wire \F_iw[31]~82_combout ;
wire \av_ld_byte3_data[7]~q ;
wire \W_rf_wr_data[31]~20_combout ;
wire \av_ld_byte3_data[6]~q ;
wire \W_rf_wr_data[30]~21_combout ;
wire \av_ld_byte3_data[5]~q ;
wire \W_rf_wr_data[29]~22_combout ;
wire \av_ld_byte3_data[4]~q ;
wire \W_rf_wr_data[28]~23_combout ;
wire \av_ld_byte3_data[3]~q ;
wire \W_rf_wr_data[27]~24_combout ;
wire \av_ld_byte3_data[2]~q ;
wire \W_rf_wr_data[26]~25_combout ;
wire \av_ld_byte3_data[1]~q ;
wire \W_rf_wr_data[25]~26_combout ;
wire \av_ld_byte3_data[0]~q ;
wire \W_rf_wr_data[24]~27_combout ;
wire \W_rf_wr_data[23]~28_combout ;
wire \W_rf_wr_data[22]~29_combout ;
wire \W_rf_wr_data[21]~30_combout ;
wire \W_rf_wr_data[20]~31_combout ;
wire \W_rf_wr_data[19]~32_combout ;
wire \W_rf_wr_data[18]~33_combout ;
wire \W_rf_wr_data[17]~34_combout ;
wire \av_ld_byte3_data_nxt~0_combout ;
wire \av_ld_byte3_data_nxt~1_combout ;
wire \av_ld_byte3_data_nxt~2_combout ;
wire \av_ld_byte3_data_nxt~3_combout ;
wire \av_ld_byte3_data_nxt~4_combout ;
wire \av_ld_byte3_data_nxt~5_combout ;
wire \av_ld_byte3_data_nxt~6_combout ;
wire \av_ld_byte3_data_nxt~7_combout ;
wire \av_ld_byte3_data_nxt~8_combout ;
wire \av_ld_byte3_data_nxt~9_combout ;
wire \av_ld_byte3_data_nxt~10_combout ;
wire \av_ld_byte3_data_nxt~11_combout ;
wire \av_ld_byte3_data_nxt~12_combout ;
wire \av_ld_byte3_data_nxt~13_combout ;
wire \av_ld_byte3_data_nxt~14_combout ;
wire \av_ld_byte3_data_nxt~15_combout ;
wire \Equal0~23_combout ;
wire \av_ld_byte0_data_nxt[0]~38_combout ;
wire \D_dst_regnum[1]~11_combout ;
wire \av_ld_byte0_data_nxt[3]~39_combout ;
wire \av_ld_byte0_data_nxt[4]~40_combout ;
wire \av_ld_byte0_data_nxt[5]~41_combout ;
wire \av_ld_byte0_data_nxt[6]~42_combout ;
wire \av_ld_byte0_data_nxt[7]~43_combout ;
wire \F_valid~0_combout ;
wire \D_valid~q ;
wire \R_valid~q ;
wire \E_new_inst~q ;
wire \F_iw[0]~14_combout ;
wire \D_iw[0]~q ;
wire \F_iw[4]~20_combout ;
wire \F_iw[4]~21_combout ;
wire \F_iw[4]~22_combout ;
wire \F_iw[4]~23_combout ;
wire \D_iw[4]~q ;
wire \F_iw[3]~24_combout ;
wire \F_iw[3]~25_combout ;
wire \F_iw[3]~26_combout ;
wire \D_iw[3]~q ;
wire \D_ctrl_st~0_combout ;
wire \F_iw[2]~27_combout ;
wire \F_iw[2]~28_combout ;
wire \F_iw[2]~29_combout ;
wire \F_iw[2]~30_combout ;
wire \D_iw[2]~q ;
wire \R_ctrl_st~q ;
wire \E_st_stall~combout ;
wire \F_iw[5]~31_combout ;
wire \F_iw[5]~32_combout ;
wire \F_iw[5]~33_combout ;
wire \F_iw[5]~34_combout ;
wire \D_iw[5]~q ;
wire \Equal0~9_combout ;
wire \W_valid~0_combout ;
wire \W_valid~q ;
wire \hbreak_pending_nxt~0_combout ;
wire \hbreak_pending~q ;
wire \wait_for_one_post_bret_inst~0_combout ;
wire \wait_for_one_post_bret_inst~q ;
wire \hbreak_req~0_combout ;
wire \F_iw[14]~35_combout ;
wire \F_iw[14]~36_combout ;
wire \F_iw[14]~83_combout ;
wire \D_iw[14]~q ;
wire \F_iw[15]~37_combout ;
wire \F_iw[15]~38_combout ;
wire \D_iw[15]~q ;
wire \D_op_opx_rsv63~0_combout ;
wire \F_iw[11]~39_combout ;
wire \D_iw[11]~q ;
wire \F_iw[13]~40_combout ;
wire \F_iw[13]~41_combout ;
wire \D_iw[13]~q ;
wire \F_iw[16]~42_combout ;
wire \F_iw[16]~43_combout ;
wire \D_iw[16]~q ;
wire \F_iw[12]~44_combout ;
wire \F_iw[12]~45_combout ;
wire \D_iw[12]~q ;
wire \Equal62~7_combout ;
wire \Equal62~9_combout ;
wire \Equal62~10_combout ;
wire \D_ctrl_shift_rot~0_combout ;
wire \D_ctrl_shift_logical~0_combout ;
wire \D_ctrl_shift_rot~1_combout ;
wire \Equal62~14_combout ;
wire \D_ctrl_shift_rot~2_combout ;
wire \D_ctrl_shift_rot~3_combout ;
wire \R_ctrl_shift_rot~q ;
wire \E_shift_rot_cnt[0]~5_combout ;
wire \D_ctrl_hi_imm16~0_combout ;
wire \D_ctrl_hi_imm16~1_combout ;
wire \R_ctrl_hi_imm16~q ;
wire \D_ctrl_alu_force_xor~14_combout ;
wire \Equal0~14_combout ;
wire \Equal0~15_combout ;
wire \D_ctrl_implicit_dst_eretaddr~3_combout ;
wire \Equal62~5_combout ;
wire \Equal62~12_combout ;
wire \D_ctrl_force_src2_zero~0_combout ;
wire \Equal62~3_combout ;
wire \D_ctrl_force_src2_zero~1_combout ;
wire \Equal62~4_combout ;
wire \D_ctrl_uncond_cti_non_br~1_combout ;
wire \Equal0~12_combout ;
wire \Equal62~6_combout ;
wire \D_ctrl_exception~4_combout ;
wire \Equal62~8_combout ;
wire \Equal0~5_combout ;
wire \D_op_opx_rsv17~0_combout ;
wire \D_ctrl_exception~5_combout ;
wire \Equal62~0_combout ;
wire \Equal62~2_combout ;
wire \D_op_opx_rsv00~0_combout ;
wire \D_ctrl_exception~6_combout ;
wire \D_ctrl_exception~7_combout ;
wire \D_ctrl_exception~8_combout ;
wire \D_ctrl_exception~9_combout ;
wire \D_ctrl_exception~10_combout ;
wire \Equal62~1_combout ;
wire \D_ctrl_exception~11_combout ;
wire \Equal62~11_combout ;
wire \D_ctrl_exception~12_combout ;
wire \Equal62~13_combout ;
wire \D_ctrl_exception~13_combout ;
wire \Equal0~10_combout ;
wire \D_ctrl_exception~14_combout ;
wire \D_ctrl_exception~15_combout ;
wire \Equal0~11_combout ;
wire \Equal0~7_combout ;
wire \D_ctrl_jmp_direct~0_combout ;
wire \D_ctrl_retaddr~0_combout ;
wire \D_ctrl_retaddr~1_combout ;
wire \D_ctrl_retaddr~2_combout ;
wire \D_ctrl_force_src2_zero~2_combout ;
wire \Equal0~21_combout ;
wire \D_ctrl_force_src2_zero~3_combout ;
wire \D_ctrl_force_src2_zero~4_combout ;
wire \D_ctrl_force_src2_zero~5_combout ;
wire \D_ctrl_force_src2_zero~6_combout ;
wire \R_ctrl_force_src2_zero~q ;
wire \R_src2_lo[4]~3_combout ;
wire \F_iw[6]~58_combout ;
wire \F_iw[6]~59_combout ;
wire \F_iw[6]~60_combout ;
wire \F_iw[6]~61_combout ;
wire \D_iw[6]~q ;
wire \D_ctrl_implicit_dst_eretaddr~0_combout ;
wire \D_ctrl_unsigned_lo_imm16~2_combout ;
wire \D_ctrl_unsigned_lo_imm16~5_combout ;
wire \D_ctrl_b_is_dst~0_combout ;
wire \D_ctrl_b_is_dst~1_combout ;
wire \D_ctrl_b_is_dst~2_combout ;
wire \Equal0~18_combout ;
wire \R_src2_use_imm~0_combout ;
wire \R_ctrl_br_nxt~0_combout ;
wire \R_ctrl_br_nxt~1_combout ;
wire \R_src2_use_imm~1_combout ;
wire \R_src2_use_imm~q ;
wire \D_ctrl_src_imm5_shift_rot~0_combout ;
wire \D_ctrl_src_imm5_shift_rot~1_combout ;
wire \R_ctrl_src_imm5_shift_rot~q ;
wire \R_src2_lo~4_combout ;
wire \R_src2_lo[0]~9_combout ;
wire \E_src2[0]~q ;
wire \E_shift_rot_cnt[0]~q ;
wire \E_shift_rot_cnt[0]~6 ;
wire \E_shift_rot_cnt[1]~7_combout ;
wire \F_iw[7]~54_combout ;
wire \F_iw[7]~55_combout ;
wire \F_iw[7]~56_combout ;
wire \F_iw[7]~57_combout ;
wire \D_iw[7]~q ;
wire \R_src2_lo[1]~8_combout ;
wire \E_src2[1]~q ;
wire \E_shift_rot_cnt[1]~q ;
wire \E_shift_rot_cnt[1]~8 ;
wire \E_shift_rot_cnt[2]~9_combout ;
wire \F_iw[8]~51_combout ;
wire \F_iw[8]~52_combout ;
wire \F_iw[8]~53_combout ;
wire \D_iw[8]~q ;
wire \R_src2_lo[2]~7_combout ;
wire \E_src2[2]~q ;
wire \E_shift_rot_cnt[2]~q ;
wire \E_stall~0_combout ;
wire \E_shift_rot_cnt[2]~10 ;
wire \E_shift_rot_cnt[3]~11_combout ;
wire \F_iw[9]~48_combout ;
wire \F_iw[9]~49_combout ;
wire \F_iw[9]~50_combout ;
wire \D_iw[9]~q ;
wire \R_src2_lo[3]~6_combout ;
wire \E_src2[3]~q ;
wire \E_shift_rot_cnt[3]~q ;
wire \E_shift_rot_cnt[3]~12 ;
wire \E_shift_rot_cnt[4]~13_combout ;
wire \F_iw[10]~46_combout ;
wire \F_iw[10]~47_combout ;
wire \D_iw[10]~q ;
wire \R_src2_lo[4]~5_combout ;
wire \E_src2[4]~q ;
wire \E_shift_rot_cnt[4]~q ;
wire \E_stall~1_combout ;
wire \E_stall~2_combout ;
wire \D_ctrl_ld_signed~0_combout ;
wire \D_ctrl_ld~2_combout ;
wire \D_ctrl_ld~3_combout ;
wire \R_ctrl_ld~q ;
wire \av_ld_waiting_for_data~q ;
wire \av_ld_aligning_data_nxt~0_combout ;
wire \av_ld_waiting_for_data_nxt~0_combout ;
wire \D_ctrl_mem16~0_combout ;
wire \av_ld_align_cycle_nxt[0]~0_combout ;
wire \av_ld_align_cycle[0]~q ;
wire \av_ld_align_cycle_nxt[1]~1_combout ;
wire \av_ld_align_cycle[1]~q ;
wire \av_ld_aligning_data_nxt~1_combout ;
wire \av_ld_aligning_data~q ;
wire \D_ctrl_mem32~0_combout ;
wire \av_ld_aligning_data_nxt~2_combout ;
wire \E_stall~3_combout ;
wire \E_stall~4_combout ;
wire \E_valid_from_R~0_combout ;
wire \E_valid_from_R~q ;
wire \D_ctrl_jmp_direct~1_combout ;
wire \R_ctrl_jmp_direct~q ;
wire \R_ctrl_br~q ;
wire \D_ctrl_retaddr~3_combout ;
wire \D_ctrl_retaddr~4_combout ;
wire \D_ctrl_retaddr~5_combout ;
wire \Equal0~13_combout ;
wire \D_ctrl_retaddr~6_combout ;
wire \D_ctrl_retaddr~7_combout ;
wire \D_ctrl_retaddr~8_combout ;
wire \R_ctrl_retaddr~q ;
wire \R_src1~35_combout ;
wire \R_src1[0]~37_combout ;
wire \E_src1[0]~q ;
wire \Equal135~0_combout ;
wire \Equal135~1_combout ;
wire \D_op_wrctl~combout ;
wire \R_ctrl_wrctl_inst~q ;
wire \W_ienable_reg_nxt~0_combout ;
wire \W_ienable_reg[0]~q ;
wire \W_ipending_reg_nxt[0]~0_combout ;
wire \W_ipending_reg[0]~q ;
wire \R_src1[1]~36_combout ;
wire \E_src1[1]~q ;
wire \W_ienable_reg[1]~q ;
wire \W_ipending_reg_nxt[1]~1_combout ;
wire \W_ipending_reg[1]~q ;
wire \E_wrctl_status~1_combout ;
wire \E_wrctl_estatus~0_combout ;
wire \D_ctrl_exception~0_combout ;
wire \D_ctrl_exception~1_combout ;
wire \D_ctrl_exception~2_combout ;
wire \D_ctrl_exception~3_combout ;
wire \D_ctrl_implicit_dst_eretaddr~1_combout ;
wire \D_ctrl_implicit_dst_eretaddr~2_combout ;
wire \D_ctrl_implicit_dst_eretaddr~4_combout ;
wire \D_ctrl_exception~16_combout ;
wire \R_ctrl_exception~q ;
wire \W_estatus_reg_inst_nxt~0_combout ;
wire \W_estatus_reg_inst_nxt~1_combout ;
wire \W_estatus_reg~q ;
wire \E_wrctl_bstatus~0_combout ;
wire \W_bstatus_reg_inst_nxt~0_combout ;
wire \D_ctrl_break~0_combout ;
wire \R_ctrl_break~q ;
wire \W_bstatus_reg_inst_nxt~1_combout ;
wire \W_bstatus_reg~q ;
wire \E_wrctl_status~0_combout ;
wire \W_status_reg_pie_inst_nxt~0_combout ;
wire \W_status_reg_pie_inst_nxt~1_combout ;
wire \D_op_eret~combout ;
wire \F_pc_sel_nxt.10~1_combout ;
wire \W_status_reg_pie_inst_nxt~2_combout ;
wire \W_status_reg_pie~q ;
wire \D_iw[26]~0_combout ;
wire \D_iw[26]~1_combout ;
wire \F_iw[1]~15_combout ;
wire \F_iw[1]~16_combout ;
wire \F_iw[1]~17_combout ;
wire \F_iw[1]~18_combout ;
wire \F_iw[1]~19_combout ;
wire \D_iw[1]~q ;
wire \Equal0~4_combout ;
wire \D_op_cmpge~0_combout ;
wire \Equal0~6_combout ;
wire \D_ctrl_alu_subtract~2_combout ;
wire \D_ctrl_alu_subtract~3_combout ;
wire \D_ctrl_alu_subtract~4_combout ;
wire \D_ctrl_alu_subtract~5_combout ;
wire \E_alu_sub~0_combout ;
wire \E_alu_sub~q ;
wire \E_src2[13]~15_combout ;
wire \R_src2_lo[7]~0_combout ;
wire \E_src2[7]~q ;
wire \Add1~0_combout ;
wire \R_src1~34_combout ;
wire \E_src1[7]~9_combout ;
wire \F_pc_plus_one[0]~1 ;
wire \F_pc_plus_one[1]~3 ;
wire \F_pc_plus_one[2]~5 ;
wire \F_pc_plus_one[3]~7 ;
wire \F_pc_plus_one[4]~9 ;
wire \F_pc_plus_one[5]~10_combout ;
wire \E_src1[7]~q ;
wire \R_src2_lo[6]~1_combout ;
wire \E_src2[6]~q ;
wire \Add1~1_combout ;
wire \E_src1[6]~10_combout ;
wire \F_pc_plus_one[4]~8_combout ;
wire \E_src1[6]~q ;
wire \R_src2_lo[5]~2_combout ;
wire \E_src2[5]~q ;
wire \Add1~2_combout ;
wire \E_src1[5]~11_combout ;
wire \F_pc_plus_one[3]~6_combout ;
wire \E_src1[5]~q ;
wire \Add1~3_combout ;
wire \E_src1[4]~12_combout ;
wire \F_pc_plus_one[2]~4_combout ;
wire \E_src1[4]~q ;
wire \Add1~4_combout ;
wire \E_src1[3]~14_combout ;
wire \F_pc_plus_one[1]~2_combout ;
wire \E_src1[3]~q ;
wire \Add1~5_combout ;
wire \E_src1[2]~13_combout ;
wire \F_pc_plus_one[0]~0_combout ;
wire \E_src1[2]~q ;
wire \Add1~6_combout ;
wire \Add1~7_combout ;
wire \Add1~9_cout ;
wire \Add1~11 ;
wire \Add1~13 ;
wire \Add1~15 ;
wire \Add1~17 ;
wire \Add1~19 ;
wire \Add1~21 ;
wire \Add1~23 ;
wire \Add1~24_combout ;
wire \D_logic_op_raw[1]~0_combout ;
wire \D_ctrl_alu_force_xor~10_combout ;
wire \D_ctrl_alu_force_xor~11_combout ;
wire \D_ctrl_alu_force_xor~13_combout ;
wire \D_ctrl_alu_force_xor~12_combout ;
wire \D_logic_op[1]~0_combout ;
wire \R_logic_op[1]~q ;
wire \D_logic_op[0]~1_combout ;
wire \R_logic_op[0]~q ;
wire \E_logic_result[7]~0_combout ;
wire \Equal0~16_combout ;
wire \Equal0~17_combout ;
wire \D_ctrl_logic~0_combout ;
wire \D_ctrl_logic~combout ;
wire \R_ctrl_logic~q ;
wire \W_alu_result[7]~9_combout ;
wire \D_ctrl_shift_rot_right~0_combout ;
wire \D_ctrl_shift_rot_right~1_combout ;
wire \R_ctrl_shift_rot_right~q ;
wire \E_shift_rot_result_nxt[6]~12_combout ;
wire \E_shift_rot_result[6]~q ;
wire \E_shift_rot_result_nxt[5]~11_combout ;
wire \E_shift_rot_result[5]~q ;
wire \E_shift_rot_result_nxt[4]~10_combout ;
wire \E_shift_rot_result[4]~q ;
wire \E_shift_rot_result_nxt[3]~14_combout ;
wire \E_shift_rot_result[3]~q ;
wire \E_shift_rot_result_nxt[2]~13_combout ;
wire \E_shift_rot_result[2]~q ;
wire \E_shift_rot_result_nxt[1]~16_combout ;
wire \E_shift_rot_result[1]~q ;
wire \E_shift_rot_result_nxt[0]~17_combout ;
wire \E_shift_rot_result[0]~q ;
wire \R_ctrl_rot_right_nxt~0_combout ;
wire \R_ctrl_rot_right~q ;
wire \D_ctrl_shift_logical~1_combout ;
wire \D_ctrl_shift_logical~2_combout ;
wire \R_ctrl_shift_logical~q ;
wire \E_shift_rot_fill_bit~0_combout ;
wire \E_shift_rot_result_nxt[31]~19_combout ;
wire \R_src1[31]~38_combout ;
wire \E_src1[31]~q ;
wire \E_shift_rot_result[31]~q ;
wire \E_shift_rot_result_nxt[30]~21_combout ;
wire \R_src1[30]~39_combout ;
wire \E_src1[30]~q ;
wire \E_shift_rot_result[30]~q ;
wire \E_shift_rot_result_nxt[29]~22_combout ;
wire \R_src1[29]~40_combout ;
wire \E_src1[29]~q ;
wire \E_shift_rot_result[29]~q ;
wire \E_shift_rot_result_nxt[28]~23_combout ;
wire \R_src1[28]~41_combout ;
wire \E_src1[28]~q ;
wire \E_shift_rot_result[28]~q ;
wire \E_shift_rot_result_nxt[27]~24_combout ;
wire \R_src1[27]~42_combout ;
wire \E_src1[27]~q ;
wire \E_shift_rot_result[27]~q ;
wire \E_shift_rot_result_nxt[26]~25_combout ;
wire \R_src1[26]~43_combout ;
wire \E_src1[26]~q ;
wire \E_shift_rot_result[26]~q ;
wire \E_shift_rot_result_nxt[25]~26_combout ;
wire \R_src1[25]~44_combout ;
wire \E_src1[25]~q ;
wire \E_shift_rot_result[25]~q ;
wire \E_shift_rot_result_nxt[24]~27_combout ;
wire \R_src1[24]~45_combout ;
wire \E_src1[24]~q ;
wire \E_shift_rot_result[24]~q ;
wire \E_shift_rot_result_nxt[23]~28_combout ;
wire \R_src1[23]~46_combout ;
wire \E_src1[23]~q ;
wire \E_shift_rot_result[23]~q ;
wire \E_shift_rot_result_nxt[22]~29_combout ;
wire \R_src1[22]~47_combout ;
wire \E_src1[22]~q ;
wire \E_shift_rot_result[22]~q ;
wire \E_shift_rot_result_nxt[21]~30_combout ;
wire \R_src1[21]~48_combout ;
wire \E_src1[21]~q ;
wire \E_shift_rot_result[21]~q ;
wire \E_shift_rot_result_nxt[20]~31_combout ;
wire \R_src1[20]~49_combout ;
wire \E_src1[20]~q ;
wire \E_shift_rot_result[20]~q ;
wire \E_shift_rot_result_nxt[19]~20_combout ;
wire \R_src1[19]~50_combout ;
wire \E_src1[19]~q ;
wire \E_shift_rot_result[19]~q ;
wire \E_shift_rot_result_nxt[18]~18_combout ;
wire \R_src1[18]~51_combout ;
wire \E_src1[18]~q ;
wire \E_shift_rot_result[18]~q ;
wire \E_shift_rot_result_nxt[17]~15_combout ;
wire \R_src1[17]~52_combout ;
wire \E_src1[17]~q ;
wire \E_shift_rot_result[17]~q ;
wire \E_shift_rot_result_nxt[16]~1_combout ;
wire \F_iw[20]~64_combout ;
wire \F_iw[20]~65_combout ;
wire \D_iw[20]~q ;
wire \E_src1[16]~0_combout ;
wire \F_pc_plus_one[5]~11 ;
wire \F_pc_plus_one[6]~13 ;
wire \F_pc_plus_one[7]~15 ;
wire \F_pc_plus_one[8]~17 ;
wire \F_pc_plus_one[9]~19 ;
wire \F_pc_plus_one[10]~21 ;
wire \F_pc_plus_one[11]~23 ;
wire \F_pc_plus_one[12]~25 ;
wire \F_pc_plus_one[13]~27 ;
wire \F_pc_plus_one[14]~28_combout ;
wire \E_src1[16]~q ;
wire \E_shift_rot_result[16]~q ;
wire \E_shift_rot_result_nxt[15]~2_combout ;
wire \F_iw[19]~66_combout ;
wire \F_iw[19]~67_combout ;
wire \D_iw[19]~q ;
wire \E_src1[15]~1_combout ;
wire \F_pc_plus_one[13]~26_combout ;
wire \E_src1[15]~q ;
wire \E_shift_rot_result[15]~q ;
wire \E_shift_rot_result_nxt[14]~3_combout ;
wire \F_iw[18]~68_combout ;
wire \F_iw[18]~69_combout ;
wire \F_iw[18]~70_combout ;
wire \D_iw[18]~q ;
wire \E_src1[14]~2_combout ;
wire \F_pc_plus_one[12]~24_combout ;
wire \E_src1[14]~q ;
wire \E_shift_rot_result[14]~q ;
wire \E_shift_rot_result_nxt[13]~4_combout ;
wire \F_iw[17]~71_combout ;
wire \F_iw[17]~72_combout ;
wire \F_iw[17]~84_combout ;
wire \D_iw[17]~q ;
wire \E_src1[13]~3_combout ;
wire \F_pc_plus_one[11]~22_combout ;
wire \E_src1[13]~q ;
wire \E_shift_rot_result[13]~q ;
wire \E_shift_rot_result_nxt[12]~5_combout ;
wire \E_src1[12]~4_combout ;
wire \F_pc_plus_one[10]~20_combout ;
wire \E_src1[12]~q ;
wire \E_shift_rot_result[12]~q ;
wire \E_shift_rot_result_nxt[11]~6_combout ;
wire \E_src1[11]~5_combout ;
wire \F_pc_plus_one[9]~18_combout ;
wire \E_src1[11]~q ;
wire \E_shift_rot_result[11]~q ;
wire \E_shift_rot_result_nxt[10]~7_combout ;
wire \E_src1[10]~6_combout ;
wire \F_pc_plus_one[8]~16_combout ;
wire \E_src1[10]~q ;
wire \E_shift_rot_result[10]~q ;
wire \E_shift_rot_result_nxt[9]~8_combout ;
wire \E_src1[9]~7_combout ;
wire \F_pc_plus_one[7]~14_combout ;
wire \E_src1[9]~q ;
wire \E_shift_rot_result[9]~q ;
wire \E_shift_rot_result_nxt[8]~9_combout ;
wire \E_src1[8]~8_combout ;
wire \F_pc_plus_one[6]~12_combout ;
wire \E_src1[8]~q ;
wire \E_shift_rot_result[8]~q ;
wire \E_shift_rot_result_nxt[7]~0_combout ;
wire \E_shift_rot_result[7]~q ;
wire \D_op_rdctl~combout ;
wire \R_ctrl_rd_ctl_reg~q ;
wire \Equal0~8_combout ;
wire \D_ctrl_br_cmp~2_combout ;
wire \D_ctrl_br_cmp~5_combout ;
wire \D_ctrl_br_cmp~3_combout ;
wire \D_ctrl_br_cmp~4_combout ;
wire \R_ctrl_br_cmp~q ;
wire \E_alu_result~0_combout ;
wire \F_iw[21]~62_combout ;
wire \F_iw[21]~63_combout ;
wire \D_iw[21]~q ;
wire \E_src2[16]~0_combout ;
wire \D_ctrl_unsigned_lo_imm16~3_combout ;
wire \D_ctrl_unsigned_lo_imm16~4_combout ;
wire \R_ctrl_unsigned_lo_imm16~q ;
wire \R_src2_hi~0_combout ;
wire \E_src2[16]~q ;
wire \Add1~26_combout ;
wire \R_src2_lo[15]~10_combout ;
wire \E_src2[15]~q ;
wire \Add1~27_combout ;
wire \R_src2_lo[14]~11_combout ;
wire \E_src2[14]~q ;
wire \Add1~28_combout ;
wire \R_src2_lo[13]~12_combout ;
wire \E_src2[13]~q ;
wire \Add1~29_combout ;
wire \R_src2_lo[12]~13_combout ;
wire \E_src2[12]~q ;
wire \Add1~30_combout ;
wire \R_src2_lo[11]~14_combout ;
wire \E_src2[11]~q ;
wire \Add1~31_combout ;
wire \R_src2_lo[10]~15_combout ;
wire \E_src2[10]~q ;
wire \Add1~32_combout ;
wire \R_src2_lo[9]~16_combout ;
wire \E_src2[9]~q ;
wire \Add1~33_combout ;
wire \R_src2_lo[8]~17_combout ;
wire \E_src2[8]~q ;
wire \Add1~34_combout ;
wire \Add1~25 ;
wire \Add1~36 ;
wire \Add1~38 ;
wire \Add1~40 ;
wire \Add1~42 ;
wire \Add1~44 ;
wire \Add1~46 ;
wire \Add1~48 ;
wire \Add1~50 ;
wire \Add1~51_combout ;
wire \E_logic_result[16]~1_combout ;
wire \W_alu_result[16]~0_combout ;
wire \Add1~49_combout ;
wire \E_logic_result[15]~2_combout ;
wire \W_alu_result[15]~1_combout ;
wire \Add1~47_combout ;
wire \E_logic_result[14]~3_combout ;
wire \W_alu_result[14]~2_combout ;
wire \Add1~45_combout ;
wire \E_logic_result[13]~4_combout ;
wire \W_alu_result[13]~3_combout ;
wire \Add1~43_combout ;
wire \E_logic_result[12]~5_combout ;
wire \W_alu_result[12]~4_combout ;
wire \Add1~41_combout ;
wire \E_logic_result[11]~6_combout ;
wire \W_alu_result[11]~5_combout ;
wire \Add1~39_combout ;
wire \E_logic_result[10]~7_combout ;
wire \W_alu_result[10]~6_combout ;
wire \Add1~37_combout ;
wire \E_logic_result[9]~8_combout ;
wire \W_alu_result[9]~7_combout ;
wire \Add1~35_combout ;
wire \E_logic_result[8]~9_combout ;
wire \W_alu_result[8]~8_combout ;
wire \Add1~18_combout ;
wire \E_logic_result[4]~10_combout ;
wire \W_alu_result[4]~12_combout ;
wire \Add1~20_combout ;
wire \E_logic_result[5]~11_combout ;
wire \W_alu_result[5]~11_combout ;
wire \Add1~22_combout ;
wire \E_logic_result[6]~12_combout ;
wire \W_alu_result[6]~10_combout ;
wire \Add1~14_combout ;
wire \E_logic_result[2]~13_combout ;
wire \W_alu_result[2]~13_combout ;
wire \Add1~16_combout ;
wire \E_logic_result[3]~14_combout ;
wire \W_alu_result[3]~14_combout ;
wire \D_ctrl_mem16~1_combout ;
wire \d_writedata[24]~0_combout ;
wire \D_ctrl_mem8~0_combout ;
wire \D_ctrl_mem8~1_combout ;
wire \d_writedata[25]~1_combout ;
wire \d_writedata[26]~2_combout ;
wire \d_writedata[27]~3_combout ;
wire \d_writedata[28]~4_combout ;
wire \d_writedata[29]~5_combout ;
wire \d_writedata[30]~6_combout ;
wire \d_writedata[31]~7_combout ;
wire \i_read_nxt~0_combout ;
wire \D_ctrl_uncond_cti_non_br~0_combout ;
wire \D_ctrl_uncond_cti_non_br~2_combout ;
wire \R_ctrl_uncond_cti_non_br~q ;
wire \Equal0~22_combout ;
wire \R_ctrl_br_uncond~q ;
wire \R_compare_op[1]~q ;
wire \R_src2_hi[15]~1_combout ;
wire \R_src2_hi[15]~2_combout ;
wire \E_src2[31]~q ;
wire \E_invert_arith_src_msb~0_combout ;
wire \E_invert_arith_src_msb~1_combout ;
wire \E_invert_arith_src_msb~q ;
wire \Add1~53_combout ;
wire \E_arith_src1[31]~combout ;
wire \E_src2[30]~1_combout ;
wire \E_src2[30]~q ;
wire \Add1~54_combout ;
wire \E_src2[29]~14_combout ;
wire \E_src2[29]~q ;
wire \Add1~55_combout ;
wire \E_src2[28]~2_combout ;
wire \E_src2[28]~q ;
wire \Add1~56_combout ;
wire \E_src2[27]~3_combout ;
wire \E_src2[27]~q ;
wire \Add1~57_combout ;
wire \E_src2[26]~4_combout ;
wire \E_src2[26]~q ;
wire \Add1~58_combout ;
wire \E_src2[25]~5_combout ;
wire \E_src2[25]~q ;
wire \Add1~59_combout ;
wire \E_src2[24]~6_combout ;
wire \E_src2[24]~q ;
wire \Add1~60_combout ;
wire \E_src2[23]~7_combout ;
wire \E_src2[23]~q ;
wire \Add1~61_combout ;
wire \E_src2[22]~8_combout ;
wire \E_src2[22]~q ;
wire \Add1~62_combout ;
wire \E_src2[21]~9_combout ;
wire \E_src2[21]~q ;
wire \Add1~63_combout ;
wire \E_src2[20]~10_combout ;
wire \E_src2[20]~q ;
wire \Add1~64_combout ;
wire \E_src2[19]~11_combout ;
wire \E_src2[19]~q ;
wire \Add1~65_combout ;
wire \E_src2[18]~12_combout ;
wire \E_src2[18]~q ;
wire \Add1~66_combout ;
wire \E_src2[17]~13_combout ;
wire \E_src2[17]~q ;
wire \Add1~67_combout ;
wire \Add1~52 ;
wire \Add1~69 ;
wire \Add1~71 ;
wire \Add1~73 ;
wire \Add1~75 ;
wire \Add1~77 ;
wire \Add1~79 ;
wire \Add1~81 ;
wire \Add1~83 ;
wire \Add1~85 ;
wire \Add1~87 ;
wire \Add1~89 ;
wire \Add1~91 ;
wire \Add1~93 ;
wire \Add1~95 ;
wire \Add1~97 ;
wire \Add1~98_combout ;
wire \Equal127~0_combout ;
wire \Equal127~1_combout ;
wire \Equal127~2_combout ;
wire \Equal127~3_combout ;
wire \E_logic_result[31]~15_combout ;
wire \Equal127~4_combout ;
wire \E_logic_result[30]~16_combout ;
wire \E_logic_result[28]~17_combout ;
wire \E_logic_result[27]~18_combout ;
wire \E_logic_result[26]~19_combout ;
wire \Equal127~5_combout ;
wire \E_logic_result[25]~20_combout ;
wire \E_logic_result[24]~21_combout ;
wire \E_logic_result[23]~22_combout ;
wire \E_logic_result[22]~23_combout ;
wire \Equal127~6_combout ;
wire \E_logic_result[21]~24_combout ;
wire \E_logic_result[20]~25_combout ;
wire \E_logic_result[19]~26_combout ;
wire \E_logic_result[18]~27_combout ;
wire \Equal127~7_combout ;
wire \E_logic_result[17]~28_combout ;
wire \E_logic_result[1]~29_combout ;
wire \E_logic_result[0]~30_combout ;
wire \E_logic_result[29]~31_combout ;
wire \Equal127~8_combout ;
wire \Equal127~9_combout ;
wire \Equal127~10_combout ;
wire \D_logic_op_raw[0]~1_combout ;
wire \R_compare_op[0]~q ;
wire \E_cmp_result~0_combout ;
wire \W_cmp_result~q ;
wire \F_pc_sel_nxt~0_combout ;
wire \F_pc_sel_nxt.10~0_combout ;
wire \F_pc_no_crst_nxt[5]~0_combout ;
wire \F_pc_no_crst_nxt[14]~1_combout ;
wire \F_pc_no_crst_nxt[14]~2_combout ;
wire \F_pc_no_crst_nxt[13]~3_combout ;
wire \F_pc_no_crst_nxt[13]~4_combout ;
wire \F_pc_no_crst_nxt[12]~5_combout ;
wire \F_pc_no_crst_nxt[11]~6_combout ;
wire \F_pc_no_crst_nxt[10]~7_combout ;
wire \F_pc_no_crst_nxt[9]~8_combout ;
wire \F_pc_no_crst_nxt[9]~9_combout ;
wire \F_pc_no_crst_nxt[8]~10_combout ;
wire \F_pc_no_crst_nxt[7]~11_combout ;
wire \F_pc_no_crst_nxt[6]~12_combout ;
wire \F_pc_no_crst_nxt[2]~13_combout ;
wire \F_pc_no_crst_nxt[3]~14_combout ;
wire \F_pc_no_crst_nxt[4]~15_combout ;
wire \d_read_nxt~combout ;
wire \F_pc_no_crst_nxt[1]~16_combout ;
wire \F_pc_no_crst_nxt[0]~17_combout ;
wire \E_st_data[9]~0_combout ;
wire \hbreak_enabled~0_combout ;
wire \Add1~10_combout ;
wire \Add1~12_combout ;
wire \E_mem_byte_en[0]~0_combout ;
wire \d_byteenable[2]~0_combout ;
wire \E_st_data[22]~1_combout ;
wire \E_mem_byte_en[2]~1_combout ;
wire \E_st_data[23]~2_combout ;
wire \E_mem_byte_en[3]~2_combout ;
wire \E_st_data[14]~3_combout ;
wire \E_mem_byte_en[1]~3_combout ;
wire \E_st_data[15]~4_combout ;
wire \E_st_data[11]~5_combout ;
wire \E_st_data[13]~6_combout ;
wire \E_st_data[16]~7_combout ;
wire \E_st_data[12]~8_combout ;
wire \E_st_data[10]~9_combout ;
wire \E_st_data[8]~10_combout ;
wire \E_st_data[21]~11_combout ;
wire \E_st_data[20]~12_combout ;
wire \E_st_data[19]~13_combout ;
wire \E_st_data[18]~14_combout ;
wire \E_st_data[17]~15_combout ;


processor_processor_nios2_gen2_0_cpu_nios2_oci the_processor_nios2_gen2_0_cpu_nios2_oci(
	.sr_0(sr_0),
	.jtag_break(\the_processor_nios2_gen2_0_cpu_nios2_oci|the_processor_nios2_gen2_0_cpu_nios2_oci_debug|jtag_break~q ),
	.readdata_0(readdata_0),
	.readdata_1(readdata_1),
	.readdata_3(readdata_3),
	.readdata_2(readdata_2),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.r_sync_rst(r_sync_rst),
	.saved_grant_0(saved_grant_0),
	.waitrequest(debug_mem_slave_waitrequest),
	.mem_used_1(mem_used_1),
	.uav_write(uav_write),
	.WideOr1(WideOr15),
	.rf_source_valid(rf_source_valid),
	.hbreak_enabled(hbreak_enabled1),
	.address_nxt({src_data_46,src_data_45,src_data_44,src_data_43,src_data_42,src_data_41,src_data_40,src_data_39,src_data_38}),
	.r_early_rst(r_early_rst),
	.oci_ienable_0(\the_processor_nios2_gen2_0_cpu_nios2_oci|the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[0]~q ),
	.oci_ienable_1(\the_processor_nios2_gen2_0_cpu_nios2_oci|the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[1]~q ),
	.oci_single_step_mode(\the_processor_nios2_gen2_0_cpu_nios2_oci|the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_single_step_mode~q ),
	.readdata_22(readdata_22),
	.readdata_23(readdata_23),
	.readdata_24(readdata_24),
	.readdata_25(readdata_25),
	.readdata_26(readdata_26),
	.readdata_4(readdata_4),
	.readdata_5(readdata_5),
	.readdata_14(readdata_14),
	.readdata_15(readdata_15),
	.readdata_11(readdata_11),
	.readdata_13(readdata_13),
	.readdata_16(readdata_16),
	.readdata_12(readdata_12),
	.readdata_10(readdata_10),
	.readdata_9(readdata_9),
	.readdata_8(readdata_8),
	.readdata_7(readdata_7),
	.readdata_6(readdata_6),
	.readdata_21(readdata_21),
	.readdata_20(readdata_20),
	.readdata_19(readdata_19),
	.readdata_18(readdata_18),
	.readdata_17(readdata_17),
	.debugaccess_nxt(src_payload11),
	.writedata_nxt({src_payload50,src_payload49,src_payload48,src_payload47,src_payload46,src_payload27,src_payload26,src_payload25,src_payload24,src_payload23,src_payload41,src_payload42,src_payload43,src_payload44,src_payload45,src_payload34,src_payload31,src_payload30,src_payload33,
src_payload35,src_payload32,src_payload36,src_payload37,src_payload38,src_payload39,src_payload40,src_payload29,src_payload28,src_payload21,src_payload22,src_payload20,src_payload12}),
	.byteenable_nxt({src_data_35,src_data_34,src_data_33,src_data_32}),
	.readdata_27(readdata_27),
	.readdata_28(readdata_28),
	.readdata_29(readdata_29),
	.readdata_30(readdata_30),
	.readdata_31(readdata_31),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_1(state_1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2),
	.clk_clk(clk_clk));

processor_processor_nios2_gen2_0_cpu_register_bank_b_module processor_nios2_gen2_0_cpu_register_bank_b(
	.q_b_0(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_1(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_2(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_3(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_4(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_5(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_6(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_7(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_16(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_15(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_14(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.q_b_13(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_12(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_11(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_10(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_9(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_8(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_31(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.q_b_30(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.q_b_29(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.q_b_28(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.q_b_27(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.q_b_26(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.q_b_25(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.q_b_24(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.q_b_23(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_22(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_21(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.q_b_20(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ),
	.q_b_19(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ),
	.q_b_18(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_17(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.W_rf_wren(\W_rf_wren~combout ),
	.W_rf_wr_data_0(\W_rf_wr_data[0]~2_combout ),
	.R_dst_regnum_0(\R_dst_regnum[0]~q ),
	.R_dst_regnum_1(\R_dst_regnum[1]~q ),
	.R_dst_regnum_2(\R_dst_regnum[2]~q ),
	.R_dst_regnum_3(\R_dst_regnum[3]~q ),
	.R_dst_regnum_4(\R_dst_regnum[4]~q ),
	.D_iw_22(\D_iw[22]~q ),
	.D_iw_23(\D_iw[23]~q ),
	.D_iw_24(\D_iw[24]~q ),
	.D_iw_25(\D_iw[25]~q ),
	.D_iw_26(\D_iw[26]~q ),
	.W_rf_wr_data_1(\W_rf_wr_data[1]~4_combout ),
	.W_rf_wr_data_2(\W_rf_wr_data[2]~5_combout ),
	.W_rf_wr_data_3(\W_rf_wr_data[3]~6_combout ),
	.W_rf_wr_data_4(\W_rf_wr_data[4]~7_combout ),
	.W_rf_wr_data_5(\W_rf_wr_data[5]~8_combout ),
	.W_rf_wr_data_6(\W_rf_wr_data[6]~9_combout ),
	.W_rf_wr_data_7(\W_rf_wr_data[7]~10_combout ),
	.W_rf_wr_data_16(\W_rf_wr_data[16]~11_combout ),
	.W_rf_wr_data_15(\W_rf_wr_data[15]~12_combout ),
	.W_rf_wr_data_14(\W_rf_wr_data[14]~13_combout ),
	.W_rf_wr_data_13(\W_rf_wr_data[13]~14_combout ),
	.W_rf_wr_data_12(\W_rf_wr_data[12]~15_combout ),
	.W_rf_wr_data_11(\W_rf_wr_data[11]~16_combout ),
	.W_rf_wr_data_10(\W_rf_wr_data[10]~17_combout ),
	.W_rf_wr_data_9(\W_rf_wr_data[9]~18_combout ),
	.W_rf_wr_data_8(\W_rf_wr_data[8]~19_combout ),
	.W_rf_wr_data_31(\W_rf_wr_data[31]~20_combout ),
	.W_rf_wr_data_30(\W_rf_wr_data[30]~21_combout ),
	.W_rf_wr_data_29(\W_rf_wr_data[29]~22_combout ),
	.W_rf_wr_data_28(\W_rf_wr_data[28]~23_combout ),
	.W_rf_wr_data_27(\W_rf_wr_data[27]~24_combout ),
	.W_rf_wr_data_26(\W_rf_wr_data[26]~25_combout ),
	.W_rf_wr_data_25(\W_rf_wr_data[25]~26_combout ),
	.W_rf_wr_data_24(\W_rf_wr_data[24]~27_combout ),
	.W_rf_wr_data_23(\W_rf_wr_data[23]~28_combout ),
	.W_rf_wr_data_22(\W_rf_wr_data[22]~29_combout ),
	.W_rf_wr_data_21(\W_rf_wr_data[21]~30_combout ),
	.W_rf_wr_data_20(\W_rf_wr_data[20]~31_combout ),
	.W_rf_wr_data_19(\W_rf_wr_data[19]~32_combout ),
	.W_rf_wr_data_18(\W_rf_wr_data[18]~33_combout ),
	.W_rf_wr_data_17(\W_rf_wr_data[17]~34_combout ),
	.clk_clk(clk_clk));

processor_processor_nios2_gen2_0_cpu_register_bank_a_module processor_nios2_gen2_0_cpu_register_bank_a(
	.q_b_7(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_6(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_5(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_4(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_3(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_2(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_1(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_0(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_16(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_15(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_14(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[14] ),
	.q_b_13(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_12(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_11(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_10(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_9(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_8(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_31(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[31] ),
	.q_b_30(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[30] ),
	.q_b_29(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[29] ),
	.q_b_28(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[28] ),
	.q_b_27(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[27] ),
	.q_b_26(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[26] ),
	.q_b_25(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[25] ),
	.q_b_24(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[24] ),
	.q_b_23(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_22(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_21(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[21] ),
	.q_b_20(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[20] ),
	.q_b_19(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[19] ),
	.q_b_18(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_17(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[17] ),
	.W_rf_wren(\W_rf_wren~combout ),
	.W_rf_wr_data_0(\W_rf_wr_data[0]~2_combout ),
	.R_dst_regnum_0(\R_dst_regnum[0]~q ),
	.R_dst_regnum_1(\R_dst_regnum[1]~q ),
	.R_dst_regnum_2(\R_dst_regnum[2]~q ),
	.R_dst_regnum_3(\R_dst_regnum[3]~q ),
	.R_dst_regnum_4(\R_dst_regnum[4]~q ),
	.W_rf_wr_data_1(\W_rf_wr_data[1]~4_combout ),
	.W_rf_wr_data_2(\W_rf_wr_data[2]~5_combout ),
	.W_rf_wr_data_3(\W_rf_wr_data[3]~6_combout ),
	.W_rf_wr_data_4(\W_rf_wr_data[4]~7_combout ),
	.W_rf_wr_data_5(\W_rf_wr_data[5]~8_combout ),
	.W_rf_wr_data_6(\W_rf_wr_data[6]~9_combout ),
	.W_rf_wr_data_7(\W_rf_wr_data[7]~10_combout ),
	.D_iw_27(\D_iw[27]~q ),
	.D_iw_28(\D_iw[28]~q ),
	.D_iw_29(\D_iw[29]~q ),
	.D_iw_30(\D_iw[30]~q ),
	.D_iw_31(\D_iw[31]~q ),
	.W_rf_wr_data_16(\W_rf_wr_data[16]~11_combout ),
	.W_rf_wr_data_15(\W_rf_wr_data[15]~12_combout ),
	.W_rf_wr_data_14(\W_rf_wr_data[14]~13_combout ),
	.W_rf_wr_data_13(\W_rf_wr_data[13]~14_combout ),
	.W_rf_wr_data_12(\W_rf_wr_data[12]~15_combout ),
	.W_rf_wr_data_11(\W_rf_wr_data[11]~16_combout ),
	.W_rf_wr_data_10(\W_rf_wr_data[10]~17_combout ),
	.W_rf_wr_data_9(\W_rf_wr_data[9]~18_combout ),
	.W_rf_wr_data_8(\W_rf_wr_data[8]~19_combout ),
	.W_rf_wr_data_31(\W_rf_wr_data[31]~20_combout ),
	.W_rf_wr_data_30(\W_rf_wr_data[30]~21_combout ),
	.W_rf_wr_data_29(\W_rf_wr_data[29]~22_combout ),
	.W_rf_wr_data_28(\W_rf_wr_data[28]~23_combout ),
	.W_rf_wr_data_27(\W_rf_wr_data[27]~24_combout ),
	.W_rf_wr_data_26(\W_rf_wr_data[26]~25_combout ),
	.W_rf_wr_data_25(\W_rf_wr_data[25]~26_combout ),
	.W_rf_wr_data_24(\W_rf_wr_data[24]~27_combout ),
	.W_rf_wr_data_23(\W_rf_wr_data[23]~28_combout ),
	.W_rf_wr_data_22(\W_rf_wr_data[22]~29_combout ),
	.W_rf_wr_data_21(\W_rf_wr_data[21]~30_combout ),
	.W_rf_wr_data_20(\W_rf_wr_data[20]~31_combout ),
	.W_rf_wr_data_19(\W_rf_wr_data[19]~32_combout ),
	.W_rf_wr_data_18(\W_rf_wr_data[18]~33_combout ),
	.W_rf_wr_data_17(\W_rf_wr_data[17]~34_combout ),
	.clk_clk(clk_clk));

dffeas \W_alu_result[0] (
	.clk(clk_clk),
	.d(\W_alu_result[0]~15_combout ),
	.asdata(\E_shift_rot_result[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[0]~q ),
	.prn(vcc));
defparam \W_alu_result[0] .is_wysiwyg = "true";
defparam \W_alu_result[0] .power_up = "low";

cyclone10lp_lcell_comb \Add1~68 (
	.dataa(\Add1~67_combout ),
	.datab(\E_src1[17]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~52 ),
	.combout(\Add1~68_combout ),
	.cout(\Add1~69 ));
defparam \Add1~68 .lut_mask = 16'h96EF;
defparam \Add1~68 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add1~70 (
	.dataa(\Add1~66_combout ),
	.datab(\E_src1[18]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~69 ),
	.combout(\Add1~70_combout ),
	.cout(\Add1~71 ));
defparam \Add1~70 .lut_mask = 16'h967F;
defparam \Add1~70 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add1~72 (
	.dataa(\Add1~65_combout ),
	.datab(\E_src1[19]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~71 ),
	.combout(\Add1~72_combout ),
	.cout(\Add1~73 ));
defparam \Add1~72 .lut_mask = 16'h96EF;
defparam \Add1~72 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add1~74 (
	.dataa(\Add1~64_combout ),
	.datab(\E_src1[20]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~73 ),
	.combout(\Add1~74_combout ),
	.cout(\Add1~75 ));
defparam \Add1~74 .lut_mask = 16'h967F;
defparam \Add1~74 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add1~76 (
	.dataa(\Add1~63_combout ),
	.datab(\E_src1[21]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~75 ),
	.combout(\Add1~76_combout ),
	.cout(\Add1~77 ));
defparam \Add1~76 .lut_mask = 16'h96EF;
defparam \Add1~76 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add1~78 (
	.dataa(\Add1~62_combout ),
	.datab(\E_src1[22]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~77 ),
	.combout(\Add1~78_combout ),
	.cout(\Add1~79 ));
defparam \Add1~78 .lut_mask = 16'h967F;
defparam \Add1~78 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add1~80 (
	.dataa(\Add1~61_combout ),
	.datab(\E_src1[23]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~79 ),
	.combout(\Add1~80_combout ),
	.cout(\Add1~81 ));
defparam \Add1~80 .lut_mask = 16'h96EF;
defparam \Add1~80 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add1~82 (
	.dataa(\Add1~60_combout ),
	.datab(\E_src1[24]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~81 ),
	.combout(\Add1~82_combout ),
	.cout(\Add1~83 ));
defparam \Add1~82 .lut_mask = 16'h967F;
defparam \Add1~82 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add1~84 (
	.dataa(\Add1~59_combout ),
	.datab(\E_src1[25]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~83 ),
	.combout(\Add1~84_combout ),
	.cout(\Add1~85 ));
defparam \Add1~84 .lut_mask = 16'h96EF;
defparam \Add1~84 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add1~86 (
	.dataa(\Add1~58_combout ),
	.datab(\E_src1[26]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~85 ),
	.combout(\Add1~86_combout ),
	.cout(\Add1~87 ));
defparam \Add1~86 .lut_mask = 16'h967F;
defparam \Add1~86 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add1~88 (
	.dataa(\Add1~57_combout ),
	.datab(\E_src1[27]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~87 ),
	.combout(\Add1~88_combout ),
	.cout(\Add1~89 ));
defparam \Add1~88 .lut_mask = 16'h96EF;
defparam \Add1~88 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add1~90 (
	.dataa(\Add1~56_combout ),
	.datab(\E_src1[28]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~89 ),
	.combout(\Add1~90_combout ),
	.cout(\Add1~91 ));
defparam \Add1~90 .lut_mask = 16'h967F;
defparam \Add1~90 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add1~92 (
	.dataa(\Add1~55_combout ),
	.datab(\E_src1[29]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~91 ),
	.combout(\Add1~92_combout ),
	.cout(\Add1~93 ));
defparam \Add1~92 .lut_mask = 16'h96EF;
defparam \Add1~92 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add1~94 (
	.dataa(\Add1~54_combout ),
	.datab(\E_src1[30]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~93 ),
	.combout(\Add1~94_combout ),
	.cout(\Add1~95 ));
defparam \Add1~94 .lut_mask = 16'h967F;
defparam \Add1~94 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add1~96 (
	.dataa(\Add1~53_combout ),
	.datab(\E_arith_src1[31]~combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~95 ),
	.combout(\Add1~96_combout ),
	.cout(\Add1~97 ));
defparam \Add1~96 .lut_mask = 16'h96EF;
defparam \Add1~96 .sum_lutc_input = "cin";

dffeas \W_alu_result[1] (
	.clk(clk_clk),
	.d(\W_alu_result[1]~16_combout ),
	.asdata(\E_shift_rot_result[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[1]~q ),
	.prn(vcc));
defparam \W_alu_result[1] .is_wysiwyg = "true";
defparam \W_alu_result[1] .power_up = "low";

dffeas \av_ld_byte1_data[0] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[0]~0_combout ),
	.asdata(\av_ld_byte2_data[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[0]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[0] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[0] .power_up = "low";

cyclone10lp_lcell_comb \W_alu_result[0]~15 (
	.dataa(\Add1~10_combout ),
	.datab(\E_logic_result[0]~30_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[0]~15_combout ),
	.cout());
defparam \W_alu_result[0]~15 .lut_mask = 16'hAACC;
defparam \W_alu_result[0]~15 .sum_lutc_input = "datac";

dffeas \av_ld_byte2_data[0] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[0]~0_combout ),
	.asdata(\av_ld_byte3_data[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[0]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[0] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[0] .power_up = "low";

dffeas \av_ld_byte1_data[7] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[7]~1_combout ),
	.asdata(\av_ld_byte2_data[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[7]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[7] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[7] .power_up = "low";

dffeas \av_ld_byte1_data[6] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[6]~2_combout ),
	.asdata(\av_ld_byte2_data[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[6]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[6] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[6] .power_up = "low";

dffeas \av_ld_byte1_data[5] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[5]~3_combout ),
	.asdata(\av_ld_byte2_data[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[5]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[5] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[5] .power_up = "low";

dffeas \av_ld_byte1_data[4] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[4]~4_combout ),
	.asdata(\av_ld_byte2_data[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[4]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[4] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[4] .power_up = "low";

dffeas \av_ld_byte1_data[3] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[3]~5_combout ),
	.asdata(\av_ld_byte2_data[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[3]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[3] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[3] .power_up = "low";

dffeas \av_ld_byte1_data[2] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[2]~6_combout ),
	.asdata(\av_ld_byte2_data[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[2]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[2] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[2] .power_up = "low";

dffeas \av_ld_byte1_data[1] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[1]~7_combout ),
	.asdata(\av_ld_byte2_data[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[1]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[1] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[1] .power_up = "low";

cyclone10lp_lcell_comb \W_alu_result[1]~16 (
	.dataa(\Add1~12_combout ),
	.datab(\E_logic_result[1]~29_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[1]~16_combout ),
	.cout());
defparam \W_alu_result[1]~16 .lut_mask = 16'hAACC;
defparam \W_alu_result[1]~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte1_data[0]~0 (
	.dataa(src_data_8),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[0]~0_combout ),
	.cout());
defparam \av_ld_byte1_data[0]~0 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[0]~0 .sum_lutc_input = "datac";

dffeas \W_alu_result[31] (
	.clk(clk_clk),
	.d(\W_alu_result[31]~17_combout ),
	.asdata(\E_shift_rot_result[31]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[31]~q ),
	.prn(vcc));
defparam \W_alu_result[31] .is_wysiwyg = "true";
defparam \W_alu_result[31] .power_up = "low";

dffeas \W_alu_result[30] (
	.clk(clk_clk),
	.d(\W_alu_result[30]~18_combout ),
	.asdata(\E_shift_rot_result[30]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[30]~q ),
	.prn(vcc));
defparam \W_alu_result[30] .is_wysiwyg = "true";
defparam \W_alu_result[30] .power_up = "low";

dffeas \W_alu_result[29] (
	.clk(clk_clk),
	.d(\W_alu_result[29]~31_combout ),
	.asdata(\E_shift_rot_result[29]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[29]~q ),
	.prn(vcc));
defparam \W_alu_result[29] .is_wysiwyg = "true";
defparam \W_alu_result[29] .power_up = "low";

dffeas \W_alu_result[28] (
	.clk(clk_clk),
	.d(\W_alu_result[28]~19_combout ),
	.asdata(\E_shift_rot_result[28]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[28]~q ),
	.prn(vcc));
defparam \W_alu_result[28] .is_wysiwyg = "true";
defparam \W_alu_result[28] .power_up = "low";

dffeas \W_alu_result[27] (
	.clk(clk_clk),
	.d(\W_alu_result[27]~20_combout ),
	.asdata(\E_shift_rot_result[27]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[27]~q ),
	.prn(vcc));
defparam \W_alu_result[27] .is_wysiwyg = "true";
defparam \W_alu_result[27] .power_up = "low";

dffeas \W_alu_result[26] (
	.clk(clk_clk),
	.d(\W_alu_result[26]~21_combout ),
	.asdata(\E_shift_rot_result[26]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[26]~q ),
	.prn(vcc));
defparam \W_alu_result[26] .is_wysiwyg = "true";
defparam \W_alu_result[26] .power_up = "low";

dffeas \W_alu_result[25] (
	.clk(clk_clk),
	.d(\W_alu_result[25]~22_combout ),
	.asdata(\E_shift_rot_result[25]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[25]~q ),
	.prn(vcc));
defparam \W_alu_result[25] .is_wysiwyg = "true";
defparam \W_alu_result[25] .power_up = "low";

dffeas \W_alu_result[24] (
	.clk(clk_clk),
	.d(\W_alu_result[24]~23_combout ),
	.asdata(\E_shift_rot_result[24]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[24]~q ),
	.prn(vcc));
defparam \W_alu_result[24] .is_wysiwyg = "true";
defparam \W_alu_result[24] .power_up = "low";

dffeas \av_ld_byte2_data[7] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[7]~1_combout ),
	.asdata(\av_ld_byte3_data[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[7]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[7] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[7] .power_up = "low";

dffeas \W_alu_result[23] (
	.clk(clk_clk),
	.d(\W_alu_result[23]~24_combout ),
	.asdata(\E_shift_rot_result[23]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[23]~q ),
	.prn(vcc));
defparam \W_alu_result[23] .is_wysiwyg = "true";
defparam \W_alu_result[23] .power_up = "low";

dffeas \av_ld_byte2_data[6] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[6]~2_combout ),
	.asdata(\av_ld_byte3_data[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[6]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[6] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[6] .power_up = "low";

dffeas \W_alu_result[22] (
	.clk(clk_clk),
	.d(\W_alu_result[22]~25_combout ),
	.asdata(\E_shift_rot_result[22]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[22]~q ),
	.prn(vcc));
defparam \W_alu_result[22] .is_wysiwyg = "true";
defparam \W_alu_result[22] .power_up = "low";

dffeas \av_ld_byte2_data[5] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[5]~3_combout ),
	.asdata(\av_ld_byte3_data[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[5]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[5] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[5] .power_up = "low";

dffeas \W_alu_result[21] (
	.clk(clk_clk),
	.d(\W_alu_result[21]~26_combout ),
	.asdata(\E_shift_rot_result[21]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[21]~q ),
	.prn(vcc));
defparam \W_alu_result[21] .is_wysiwyg = "true";
defparam \W_alu_result[21] .power_up = "low";

dffeas \av_ld_byte2_data[4] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[4]~4_combout ),
	.asdata(\av_ld_byte3_data[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[4]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[4] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[4] .power_up = "low";

dffeas \W_alu_result[20] (
	.clk(clk_clk),
	.d(\W_alu_result[20]~27_combout ),
	.asdata(\E_shift_rot_result[20]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[20]~q ),
	.prn(vcc));
defparam \W_alu_result[20] .is_wysiwyg = "true";
defparam \W_alu_result[20] .power_up = "low";

dffeas \av_ld_byte2_data[3] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[3]~5_combout ),
	.asdata(\av_ld_byte3_data[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[3]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[3] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[3] .power_up = "low";

dffeas \W_alu_result[19] (
	.clk(clk_clk),
	.d(\W_alu_result[19]~28_combout ),
	.asdata(\E_shift_rot_result[19]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[19]~q ),
	.prn(vcc));
defparam \W_alu_result[19] .is_wysiwyg = "true";
defparam \W_alu_result[19] .power_up = "low";

dffeas \av_ld_byte2_data[2] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[2]~6_combout ),
	.asdata(\av_ld_byte3_data[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[2]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[2] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[2] .power_up = "low";

dffeas \W_alu_result[18] (
	.clk(clk_clk),
	.d(\W_alu_result[18]~29_combout ),
	.asdata(\E_shift_rot_result[18]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[18]~q ),
	.prn(vcc));
defparam \W_alu_result[18] .is_wysiwyg = "true";
defparam \W_alu_result[18] .power_up = "low";

dffeas \av_ld_byte2_data[1] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[1]~7_combout ),
	.asdata(\av_ld_byte3_data[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[1]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[1] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[1] .power_up = "low";

dffeas \W_alu_result[17] (
	.clk(clk_clk),
	.d(\W_alu_result[17]~30_combout ),
	.asdata(\E_shift_rot_result[17]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[17]~q ),
	.prn(vcc));
defparam \W_alu_result[17] .is_wysiwyg = "true";
defparam \W_alu_result[17] .power_up = "low";

cyclone10lp_lcell_comb \av_ld_byte2_data[0]~0 (
	.dataa(src_payload4),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[0]~0_combout ),
	.cout());
defparam \av_ld_byte2_data[0]~0 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte1_data[7]~1 (
	.dataa(src_payload5),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[7]~1_combout ),
	.cout());
defparam \av_ld_byte1_data[7]~1 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[7]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte1_data[6]~2 (
	.dataa(src_payload6),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[6]~2_combout ),
	.cout());
defparam \av_ld_byte1_data[6]~2 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[6]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte1_data[5]~3 (
	.dataa(src_payload7),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[5]~3_combout ),
	.cout());
defparam \av_ld_byte1_data[5]~3 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[5]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte1_data[4]~4 (
	.dataa(src_payload8),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[4]~4_combout ),
	.cout());
defparam \av_ld_byte1_data[4]~4 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[4]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte1_data[3]~5 (
	.dataa(src_payload9),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[3]~5_combout ),
	.cout());
defparam \av_ld_byte1_data[3]~5 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[3]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte1_data[2]~6 (
	.dataa(src_payload10),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[2]~6_combout ),
	.cout());
defparam \av_ld_byte1_data[2]~6 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[2]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte1_data[1]~7 (
	.dataa(src_data_9),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[1]~7_combout ),
	.cout());
defparam \av_ld_byte1_data[1]~7 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[1]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_alu_result[31]~17 (
	.dataa(\Add1~96_combout ),
	.datab(\E_logic_result[31]~15_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[31]~17_combout ),
	.cout());
defparam \W_alu_result[31]~17 .lut_mask = 16'hAACC;
defparam \W_alu_result[31]~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_alu_result[30]~18 (
	.dataa(\Add1~94_combout ),
	.datab(\E_logic_result[30]~16_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[30]~18_combout ),
	.cout());
defparam \W_alu_result[30]~18 .lut_mask = 16'hAACC;
defparam \W_alu_result[30]~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_alu_result[29]~31 (
	.dataa(\Add1~92_combout ),
	.datab(\E_logic_result[29]~31_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[29]~31_combout ),
	.cout());
defparam \W_alu_result[29]~31 .lut_mask = 16'hAACC;
defparam \W_alu_result[29]~31 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_alu_result[28]~19 (
	.dataa(\Add1~90_combout ),
	.datab(\E_logic_result[28]~17_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[28]~19_combout ),
	.cout());
defparam \W_alu_result[28]~19 .lut_mask = 16'hAACC;
defparam \W_alu_result[28]~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_alu_result[27]~20 (
	.dataa(\Add1~88_combout ),
	.datab(\E_logic_result[27]~18_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[27]~20_combout ),
	.cout());
defparam \W_alu_result[27]~20 .lut_mask = 16'hAACC;
defparam \W_alu_result[27]~20 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_alu_result[26]~21 (
	.dataa(\Add1~86_combout ),
	.datab(\E_logic_result[26]~19_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[26]~21_combout ),
	.cout());
defparam \W_alu_result[26]~21 .lut_mask = 16'hAACC;
defparam \W_alu_result[26]~21 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_alu_result[25]~22 (
	.dataa(\Add1~84_combout ),
	.datab(\E_logic_result[25]~20_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[25]~22_combout ),
	.cout());
defparam \W_alu_result[25]~22 .lut_mask = 16'hAACC;
defparam \W_alu_result[25]~22 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_alu_result[24]~23 (
	.dataa(\Add1~82_combout ),
	.datab(\E_logic_result[24]~21_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[24]~23_combout ),
	.cout());
defparam \W_alu_result[24]~23 .lut_mask = 16'hAACC;
defparam \W_alu_result[24]~23 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte2_data[7]~1 (
	.dataa(src_payload13),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[7]~1_combout ),
	.cout());
defparam \av_ld_byte2_data[7]~1 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[7]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_alu_result[23]~24 (
	.dataa(\Add1~80_combout ),
	.datab(\E_logic_result[23]~22_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[23]~24_combout ),
	.cout());
defparam \W_alu_result[23]~24 .lut_mask = 16'hAACC;
defparam \W_alu_result[23]~24 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte2_data[6]~2 (
	.dataa(src_payload14),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[6]~2_combout ),
	.cout());
defparam \av_ld_byte2_data[6]~2 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[6]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_alu_result[22]~25 (
	.dataa(\Add1~78_combout ),
	.datab(\E_logic_result[22]~23_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[22]~25_combout ),
	.cout());
defparam \W_alu_result[22]~25 .lut_mask = 16'hAACC;
defparam \W_alu_result[22]~25 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte2_data[5]~3 (
	.dataa(src_payload15),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[5]~3_combout ),
	.cout());
defparam \av_ld_byte2_data[5]~3 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[5]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_alu_result[21]~26 (
	.dataa(\Add1~76_combout ),
	.datab(\E_logic_result[21]~24_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[21]~26_combout ),
	.cout());
defparam \W_alu_result[21]~26 .lut_mask = 16'hAACC;
defparam \W_alu_result[21]~26 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte2_data[4]~4 (
	.dataa(src_payload16),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[4]~4_combout ),
	.cout());
defparam \av_ld_byte2_data[4]~4 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[4]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_alu_result[20]~27 (
	.dataa(\Add1~74_combout ),
	.datab(\E_logic_result[20]~25_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[20]~27_combout ),
	.cout());
defparam \W_alu_result[20]~27 .lut_mask = 16'hAACC;
defparam \W_alu_result[20]~27 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte2_data[3]~5 (
	.dataa(src_payload17),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[3]~5_combout ),
	.cout());
defparam \av_ld_byte2_data[3]~5 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[3]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_alu_result[19]~28 (
	.dataa(\Add1~72_combout ),
	.datab(\E_logic_result[19]~26_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[19]~28_combout ),
	.cout());
defparam \W_alu_result[19]~28 .lut_mask = 16'hAACC;
defparam \W_alu_result[19]~28 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte2_data[2]~6 (
	.dataa(src_payload18),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[2]~6_combout ),
	.cout());
defparam \av_ld_byte2_data[2]~6 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[2]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_alu_result[18]~29 (
	.dataa(\Add1~70_combout ),
	.datab(\E_logic_result[18]~27_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[18]~29_combout ),
	.cout());
defparam \W_alu_result[18]~29 .lut_mask = 16'hAACC;
defparam \W_alu_result[18]~29 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte2_data[1]~7 (
	.dataa(src_payload19),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[1]~7_combout ),
	.cout());
defparam \av_ld_byte2_data[1]~7 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[1]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_alu_result[17]~30 (
	.dataa(\Add1~68_combout ),
	.datab(\E_logic_result[17]~28_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[17]~30_combout ),
	.cout());
defparam \W_alu_result[17]~30 .lut_mask = 16'hAACC;
defparam \W_alu_result[17]~30 .sum_lutc_input = "datac";

dffeas R_wr_dst_reg(
	.clk(clk_clk),
	.d(\D_wr_dst_reg~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_wr_dst_reg~q ),
	.prn(vcc));
defparam R_wr_dst_reg.is_wysiwyg = "true";
defparam R_wr_dst_reg.power_up = "low";

cyclone10lp_lcell_comb W_rf_wren(
	.dataa(r_sync_rst),
	.datab(\W_valid~q ),
	.datac(\R_wr_dst_reg~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\W_rf_wren~combout ),
	.cout());
defparam W_rf_wren.lut_mask = 16'hFEFE;
defparam W_rf_wren.sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[0] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[0]~38_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[7]~0_combout ),
	.q(\av_ld_byte0_data[0]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[0] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[0] .power_up = "low";

cyclone10lp_lcell_comb \W_rf_wr_data[0]~0 (
	.dataa(\W_cmp_result~q ),
	.datab(\R_ctrl_br_cmp~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\W_rf_wr_data[0]~0_combout ),
	.cout());
defparam \W_rf_wr_data[0]~0 .lut_mask = 16'hEEEE;
defparam \W_rf_wr_data[0]~0 .sum_lutc_input = "datac";

dffeas \W_control_rd_data[0] (
	.clk(clk_clk),
	.d(\E_control_rd_data[0]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_control_rd_data[0]~q ),
	.prn(vcc));
defparam \W_control_rd_data[0] .is_wysiwyg = "true";
defparam \W_control_rd_data[0] .power_up = "low";

cyclone10lp_lcell_comb \W_rf_wr_data[0]~1 (
	.dataa(\W_control_rd_data[0]~q ),
	.datab(\W_alu_result[0]~q ),
	.datac(\R_ctrl_rd_ctl_reg~q ),
	.datad(\R_ctrl_br_cmp~q ),
	.cin(gnd),
	.combout(\W_rf_wr_data[0]~1_combout ),
	.cout());
defparam \W_rf_wr_data[0]~1 .lut_mask = 16'hACFF;
defparam \W_rf_wr_data[0]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_rf_wr_data[0]~2 (
	.dataa(\av_ld_byte0_data[0]~q ),
	.datab(\W_rf_wr_data[0]~0_combout ),
	.datac(\W_rf_wr_data[0]~1_combout ),
	.datad(\R_ctrl_ld~q ),
	.cin(gnd),
	.combout(\W_rf_wr_data[0]~2_combout ),
	.cout());
defparam \W_rf_wr_data[0]~2 .lut_mask = 16'hFAFC;
defparam \W_rf_wr_data[0]~2 .sum_lutc_input = "datac";

dffeas \R_dst_regnum[0] (
	.clk(clk_clk),
	.d(\D_dst_regnum[0]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[0]~q ),
	.prn(vcc));
defparam \R_dst_regnum[0] .is_wysiwyg = "true";
defparam \R_dst_regnum[0] .power_up = "low";

dffeas \R_dst_regnum[1] (
	.clk(clk_clk),
	.d(\D_dst_regnum[1]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[1]~q ),
	.prn(vcc));
defparam \R_dst_regnum[1] .is_wysiwyg = "true";
defparam \R_dst_regnum[1] .power_up = "low";

dffeas \R_dst_regnum[2] (
	.clk(clk_clk),
	.d(\D_dst_regnum[2]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[2]~q ),
	.prn(vcc));
defparam \R_dst_regnum[2] .is_wysiwyg = "true";
defparam \R_dst_regnum[2] .power_up = "low";

dffeas \R_dst_regnum[3] (
	.clk(clk_clk),
	.d(\D_dst_regnum[3]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[3]~q ),
	.prn(vcc));
defparam \R_dst_regnum[3] .is_wysiwyg = "true";
defparam \R_dst_regnum[3] .power_up = "low";

dffeas \R_dst_regnum[4] (
	.clk(clk_clk),
	.d(\D_dst_regnum[4]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[4]~q ),
	.prn(vcc));
defparam \R_dst_regnum[4] .is_wysiwyg = "true";
defparam \R_dst_regnum[4] .power_up = "low";

dffeas \D_iw[22] (
	.clk(clk_clk),
	.d(\F_iw[22]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[22]~q ),
	.prn(vcc));
defparam \D_iw[22] .is_wysiwyg = "true";
defparam \D_iw[22] .power_up = "low";

dffeas \D_iw[23] (
	.clk(clk_clk),
	.d(\F_iw[23]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[23]~q ),
	.prn(vcc));
defparam \D_iw[23] .is_wysiwyg = "true";
defparam \D_iw[23] .power_up = "low";

dffeas \D_iw[24] (
	.clk(clk_clk),
	.d(\F_iw[24]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[24]~q ),
	.prn(vcc));
defparam \D_iw[24] .is_wysiwyg = "true";
defparam \D_iw[24] .power_up = "low";

dffeas \D_iw[25] (
	.clk(clk_clk),
	.d(\F_iw[25]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[25]~q ),
	.prn(vcc));
defparam \D_iw[25] .is_wysiwyg = "true";
defparam \D_iw[25] .power_up = "low";

dffeas \D_iw[26] (
	.clk(clk_clk),
	.d(\F_iw[26]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[26]~q ),
	.prn(vcc));
defparam \D_iw[26] .is_wysiwyg = "true";
defparam \D_iw[26] .power_up = "low";

cyclone10lp_lcell_comb \D_ctrl_ld_signed~1 (
	.dataa(\D_iw[2]~q ),
	.datab(\D_ctrl_ld_signed~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_ld_signed~1_combout ),
	.cout());
defparam \D_ctrl_ld_signed~1 .lut_mask = 16'hEEEE;
defparam \D_ctrl_ld_signed~1 .sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[1] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[1]~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[7]~0_combout ),
	.q(\av_ld_byte0_data[1]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[1] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[1] .power_up = "low";

dffeas \W_control_rd_data[1] (
	.clk(clk_clk),
	.d(\E_control_rd_data[1]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_control_rd_data[1]~q ),
	.prn(vcc));
defparam \W_control_rd_data[1] .is_wysiwyg = "true";
defparam \W_control_rd_data[1] .power_up = "low";

cyclone10lp_lcell_comb \W_rf_wr_data[1]~3 (
	.dataa(\W_control_rd_data[1]~q ),
	.datab(\W_alu_result[1]~q ),
	.datac(\R_ctrl_rd_ctl_reg~q ),
	.datad(\R_ctrl_br_cmp~q ),
	.cin(gnd),
	.combout(\W_rf_wr_data[1]~3_combout ),
	.cout());
defparam \W_rf_wr_data[1]~3 .lut_mask = 16'hACFF;
defparam \W_rf_wr_data[1]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_rf_wr_data[1]~4 (
	.dataa(\av_ld_byte0_data[1]~q ),
	.datab(\W_rf_wr_data[1]~3_combout ),
	.datac(gnd),
	.datad(\R_ctrl_ld~q ),
	.cin(gnd),
	.combout(\W_rf_wr_data[1]~4_combout ),
	.cout());
defparam \W_rf_wr_data[1]~4 .lut_mask = 16'hAACC;
defparam \W_rf_wr_data[1]~4 .sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[2] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[2]~22_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[7]~0_combout ),
	.q(\av_ld_byte0_data[2]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[2] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[2] .power_up = "low";

cyclone10lp_lcell_comb \W_rf_wr_data[2]~5 (
	.dataa(\av_ld_byte0_data[2]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_2),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[2]~5_combout ),
	.cout());
defparam \W_rf_wr_data[2]~5 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[2]~5 .sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[3] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[3]~39_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[7]~0_combout ),
	.q(\av_ld_byte0_data[3]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[3] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[3] .power_up = "low";

cyclone10lp_lcell_comb \W_rf_wr_data[3]~6 (
	.dataa(\av_ld_byte0_data[3]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_3),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[3]~6_combout ),
	.cout());
defparam \W_rf_wr_data[3]~6 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[3]~6 .sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[4] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[4]~40_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[7]~0_combout ),
	.q(\av_ld_byte0_data[4]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[4] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[4] .power_up = "low";

cyclone10lp_lcell_comb \W_rf_wr_data[4]~7 (
	.dataa(\av_ld_byte0_data[4]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_4),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[4]~7_combout ),
	.cout());
defparam \W_rf_wr_data[4]~7 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[4]~7 .sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[5] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[5]~41_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[7]~0_combout ),
	.q(\av_ld_byte0_data[5]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[5] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[5] .power_up = "low";

cyclone10lp_lcell_comb \W_rf_wr_data[5]~8 (
	.dataa(\av_ld_byte0_data[5]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_5),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[5]~8_combout ),
	.cout());
defparam \W_rf_wr_data[5]~8 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[5]~8 .sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[6] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[6]~42_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[7]~0_combout ),
	.q(\av_ld_byte0_data[6]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[6] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[6] .power_up = "low";

cyclone10lp_lcell_comb \W_rf_wr_data[6]~9 (
	.dataa(\av_ld_byte0_data[6]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_6),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[6]~9_combout ),
	.cout());
defparam \W_rf_wr_data[6]~9 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[6]~9 .sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[7] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[7]~43_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[7]~0_combout ),
	.q(\av_ld_byte0_data[7]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[7] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[7] .power_up = "low";

cyclone10lp_lcell_comb \W_rf_wr_data[7]~10 (
	.dataa(\av_ld_byte0_data[7]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_7),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[7]~10_combout ),
	.cout());
defparam \W_rf_wr_data[7]~10 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[7]~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_wr_dst_reg~0 (
	.dataa(\Equal0~15_combout ),
	.datab(\Equal0~12_combout ),
	.datac(\D_iw[5]~q ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_wr_dst_reg~0_combout ),
	.cout());
defparam \D_wr_dst_reg~0 .lut_mask = 16'hEFFF;
defparam \D_wr_dst_reg~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_wr_dst_reg~1 (
	.dataa(\R_ctrl_br_nxt~1_combout ),
	.datab(\D_wr_dst_reg~0_combout ),
	.datac(\Equal0~18_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_wr_dst_reg~1_combout ),
	.cout());
defparam \D_wr_dst_reg~1 .lut_mask = 16'hFEFE;
defparam \D_wr_dst_reg~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_implicit_dst_eretaddr~5 (
	.dataa(\Equal62~6_combout ),
	.datab(\Equal62~12_combout ),
	.datac(\D_iw[14]~q ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~5_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~5 .lut_mask = 16'hEFFE;
defparam \D_ctrl_implicit_dst_eretaddr~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_implicit_dst_eretaddr~6 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[12]~q ),
	.datac(\D_iw[13]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~6_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~6 .lut_mask = 16'hFBFF;
defparam \D_ctrl_implicit_dst_eretaddr~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_implicit_dst_eretaddr~7 (
	.dataa(\Equal0~9_combout ),
	.datab(\D_ctrl_implicit_dst_eretaddr~5_combout ),
	.datac(\D_ctrl_exception~2_combout ),
	.datad(\D_ctrl_implicit_dst_eretaddr~6_combout ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~7_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~7 .lut_mask = 16'hFFFE;
defparam \D_ctrl_implicit_dst_eretaddr~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_implicit_dst_eretaddr~8 (
	.dataa(\D_ctrl_implicit_dst_eretaddr~7_combout ),
	.datab(\D_ctrl_exception~8_combout ),
	.datac(\D_ctrl_exception~15_combout ),
	.datad(\D_ctrl_implicit_dst_eretaddr~4_combout ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~8_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~8 .lut_mask = 16'hBFFF;
defparam \D_ctrl_implicit_dst_eretaddr~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_dst_regnum[0]~2 (
	.dataa(\D_iw[4]~q ),
	.datab(\D_iw[5]~q ),
	.datac(\Equal0~7_combout ),
	.datad(\D_ctrl_implicit_dst_eretaddr~8_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[0]~2_combout ),
	.cout());
defparam \D_dst_regnum[0]~2 .lut_mask = 16'hEFFF;
defparam \D_dst_regnum[0]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_dst_regnum[1]~3 (
	.dataa(\D_iw[23]~q ),
	.datab(\D_iw[18]~q ),
	.datac(\D_ctrl_b_is_dst~2_combout ),
	.datad(\D_ctrl_implicit_dst_eretaddr~8_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[1]~3_combout ),
	.cout());
defparam \D_dst_regnum[1]~3 .lut_mask = 16'hACFF;
defparam \D_dst_regnum[1]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_dst_regnum[0]~4 (
	.dataa(\D_iw[22]~q ),
	.datab(\D_iw[17]~q ),
	.datac(gnd),
	.datad(\D_ctrl_b_is_dst~2_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[0]~4_combout ),
	.cout());
defparam \D_dst_regnum[0]~4 .lut_mask = 16'hAACC;
defparam \D_dst_regnum[0]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal0~19 (
	.dataa(\D_dst_regnum[0]~2_combout ),
	.datab(\Equal0~23_combout ),
	.datac(\D_dst_regnum[1]~3_combout ),
	.datad(\D_dst_regnum[0]~4_combout ),
	.cin(gnd),
	.combout(\Equal0~19_combout ),
	.cout());
defparam \Equal0~19 .lut_mask = 16'hBFFF;
defparam \Equal0~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_dst_regnum[3]~5 (
	.dataa(\D_iw[25]~q ),
	.datab(\D_iw[20]~q ),
	.datac(gnd),
	.datad(\D_ctrl_b_is_dst~2_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[3]~5_combout ),
	.cout());
defparam \D_dst_regnum[3]~5 .lut_mask = 16'hAACC;
defparam \D_dst_regnum[3]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_dst_regnum[4]~6 (
	.dataa(\D_iw[26]~q ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\D_ctrl_b_is_dst~2_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[4]~6_combout ),
	.cout());
defparam \D_dst_regnum[4]~6 .lut_mask = 16'hAACC;
defparam \D_dst_regnum[4]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal0~20 (
	.dataa(\Equal0~23_combout ),
	.datab(\D_ctrl_implicit_dst_eretaddr~8_combout ),
	.datac(\D_dst_regnum[3]~5_combout ),
	.datad(\D_dst_regnum[4]~6_combout ),
	.cin(gnd),
	.combout(\Equal0~20_combout ),
	.cout());
defparam \Equal0~20 .lut_mask = 16'h7FFF;
defparam \Equal0~20 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_dst_regnum[2]~7 (
	.dataa(\D_iw[24]~q ),
	.datab(\D_iw[19]~q ),
	.datac(\D_ctrl_b_is_dst~2_combout ),
	.datad(\D_dst_regnum[0]~2_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[2]~7_combout ),
	.cout());
defparam \D_dst_regnum[2]~7 .lut_mask = 16'hACFF;
defparam \D_dst_regnum[2]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_wr_dst_reg~2 (
	.dataa(\D_wr_dst_reg~1_combout ),
	.datab(\Equal0~19_combout ),
	.datac(\Equal0~20_combout ),
	.datad(\D_dst_regnum[2]~7_combout ),
	.cin(gnd),
	.combout(\D_wr_dst_reg~2_combout ),
	.cout());
defparam \D_wr_dst_reg~2 .lut_mask = 16'hFF7F;
defparam \D_wr_dst_reg~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_rshift8~0 (
	.dataa(\W_alu_result[1]~q ),
	.datab(\W_alu_result[0]~q ),
	.datac(\av_ld_align_cycle[0]~q ),
	.datad(\av_ld_align_cycle[1]~q ),
	.cin(gnd),
	.combout(\av_ld_rshift8~0_combout ),
	.cout());
defparam \av_ld_rshift8~0 .lut_mask = 16'hEFFF;
defparam \av_ld_rshift8~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_rshift8~1 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\av_ld_rshift8~1_combout ),
	.cout());
defparam \av_ld_rshift8~1 .lut_mask = 16'hEEEE;
defparam \av_ld_rshift8~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data[7]~0 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\av_ld_rshift8~0_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data[7]~0_combout ),
	.cout());
defparam \av_ld_byte0_data[7]~0 .lut_mask = 16'hFF55;
defparam \av_ld_byte0_data[7]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_control_rd_data[0]~0 (
	.dataa(\W_estatus_reg~q ),
	.datab(\W_status_reg_pie~q ),
	.datac(\D_iw[6]~q ),
	.datad(\D_iw[8]~q ),
	.cin(gnd),
	.combout(\E_control_rd_data[0]~0_combout ),
	.cout());
defparam \E_control_rd_data[0]~0 .lut_mask = 16'hACFF;
defparam \E_control_rd_data[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_control_rd_data[0]~1 (
	.dataa(\W_bstatus_reg~q ),
	.datab(\W_ipending_reg[0]~q ),
	.datac(\D_iw[8]~q ),
	.datad(\D_iw[7]~q ),
	.cin(gnd),
	.combout(\E_control_rd_data[0]~1_combout ),
	.cout());
defparam \E_control_rd_data[0]~1 .lut_mask = 16'hEFFE;
defparam \E_control_rd_data[0]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_control_rd_data[0]~2 (
	.dataa(\E_control_rd_data[0]~0_combout ),
	.datab(\E_control_rd_data[0]~1_combout ),
	.datac(\D_iw[7]~q ),
	.datad(\D_iw[6]~q ),
	.cin(gnd),
	.combout(\E_control_rd_data[0]~2_combout ),
	.cout());
defparam \E_control_rd_data[0]~2 .lut_mask = 16'hEFFF;
defparam \E_control_rd_data[0]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_control_rd_data[0]~3 (
	.dataa(\W_ienable_reg[0]~q ),
	.datab(\Equal135~0_combout ),
	.datac(\E_control_rd_data[0]~2_combout ),
	.datad(\Equal135~1_combout ),
	.cin(gnd),
	.combout(\E_control_rd_data[0]~3_combout ),
	.cout());
defparam \E_control_rd_data[0]~3 .lut_mask = 16'hFFFE;
defparam \E_control_rd_data[0]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_dst_regnum[0]~8 (
	.dataa(\Equal0~23_combout ),
	.datab(\D_ctrl_implicit_dst_eretaddr~8_combout ),
	.datac(\D_dst_regnum[0]~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_dst_regnum[0]~8_combout ),
	.cout());
defparam \D_dst_regnum[0]~8 .lut_mask = 16'hFEFE;
defparam \D_dst_regnum[0]~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_dst_regnum[3]~9 (
	.dataa(\Equal0~23_combout ),
	.datab(\D_ctrl_implicit_dst_eretaddr~8_combout ),
	.datac(\D_dst_regnum[3]~5_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_dst_regnum[3]~9_combout ),
	.cout());
defparam \D_dst_regnum[3]~9 .lut_mask = 16'hFEFE;
defparam \D_dst_regnum[3]~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_dst_regnum[4]~10 (
	.dataa(\Equal0~23_combout ),
	.datab(\D_ctrl_implicit_dst_eretaddr~8_combout ),
	.datac(\D_dst_regnum[4]~6_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_dst_regnum[4]~10_combout ),
	.cout());
defparam \D_dst_regnum[4]~10 .lut_mask = 16'hFEFE;
defparam \D_dst_regnum[4]~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[22]~4 (
	.dataa(src1_valid1),
	.datab(src1_valid2),
	.datac(q_a_22),
	.datad(av_readdata_pre_221),
	.cin(gnd),
	.combout(\F_iw[22]~4_combout ),
	.cout());
defparam \F_iw[22]~4 .lut_mask = 16'hFFFE;
defparam \F_iw[22]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[22]~5 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[22]~4_combout ),
	.datac(src1_valid),
	.datad(av_readdata_pre_22),
	.cin(gnd),
	.combout(\F_iw[22]~5_combout ),
	.cout());
defparam \F_iw[22]~5 .lut_mask = 16'hFFFE;
defparam \F_iw[22]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[23]~6 (
	.dataa(read_latency_shift_reg_0),
	.datab(mem_74_0),
	.datac(mem_56_0),
	.datad(av_readdata_pre_23),
	.cin(gnd),
	.combout(\F_iw[23]~6_combout ),
	.cout());
defparam \F_iw[23]~6 .lut_mask = 16'hFFFE;
defparam \F_iw[23]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[23]~7 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[23]~6_combout ),
	.datac(src1_valid2),
	.datad(q_a_23),
	.cin(gnd),
	.combout(\F_iw[23]~7_combout ),
	.cout());
defparam \F_iw[23]~7 .lut_mask = 16'hFFFE;
defparam \F_iw[23]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[24]~8 (
	.dataa(read_latency_shift_reg_0),
	.datab(mem_74_0),
	.datac(mem_56_0),
	.datad(av_readdata_pre_24),
	.cin(gnd),
	.combout(\F_iw[24]~8_combout ),
	.cout());
defparam \F_iw[24]~8 .lut_mask = 16'hFFFE;
defparam \F_iw[24]~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[24]~9 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[24]~8_combout ),
	.datac(src1_valid2),
	.datad(q_a_24),
	.cin(gnd),
	.combout(\F_iw[24]~9_combout ),
	.cout());
defparam \F_iw[24]~9 .lut_mask = 16'hFFFE;
defparam \F_iw[24]~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[25]~10 (
	.dataa(read_latency_shift_reg_0),
	.datab(mem_74_0),
	.datac(mem_56_0),
	.datad(av_readdata_pre_25),
	.cin(gnd),
	.combout(\F_iw[25]~10_combout ),
	.cout());
defparam \F_iw[25]~10 .lut_mask = 16'hFFFE;
defparam \F_iw[25]~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[25]~11 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[25]~10_combout ),
	.datac(src1_valid2),
	.datad(q_a_25),
	.cin(gnd),
	.combout(\F_iw[25]~11_combout ),
	.cout());
defparam \F_iw[25]~11 .lut_mask = 16'hFFFE;
defparam \F_iw[25]~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[26]~12 (
	.dataa(read_latency_shift_reg_0),
	.datab(mem_74_0),
	.datac(mem_56_0),
	.datad(av_readdata_pre_26),
	.cin(gnd),
	.combout(\F_iw[26]~12_combout ),
	.cout());
defparam \F_iw[26]~12 .lut_mask = 16'hFFFE;
defparam \F_iw[26]~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[26]~13 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[26]~12_combout ),
	.datac(src1_valid2),
	.datad(q_a_26),
	.cin(gnd),
	.combout(\F_iw[26]~13_combout ),
	.cout());
defparam \F_iw[26]~13 .lut_mask = 16'hFFFE;
defparam \F_iw[26]~13 .sum_lutc_input = "datac";

dffeas \D_iw[27] (
	.clk(clk_clk),
	.d(\F_iw[27]~74_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[27]~q ),
	.prn(vcc));
defparam \D_iw[27] .is_wysiwyg = "true";
defparam \D_iw[27] .power_up = "low";

dffeas \D_iw[28] (
	.clk(clk_clk),
	.d(\F_iw[28]~76_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[28]~q ),
	.prn(vcc));
defparam \D_iw[28] .is_wysiwyg = "true";
defparam \D_iw[28] .power_up = "low";

dffeas \D_iw[29] (
	.clk(clk_clk),
	.d(\F_iw[29]~78_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[29]~q ),
	.prn(vcc));
defparam \D_iw[29] .is_wysiwyg = "true";
defparam \D_iw[29] .power_up = "low";

dffeas \D_iw[30] (
	.clk(clk_clk),
	.d(\F_iw[30]~80_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[30]~q ),
	.prn(vcc));
defparam \D_iw[30] .is_wysiwyg = "true";
defparam \D_iw[30] .power_up = "low";

dffeas \D_iw[31] (
	.clk(clk_clk),
	.d(\F_iw[31]~82_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[31]~q ),
	.prn(vcc));
defparam \D_iw[31] .is_wysiwyg = "true";
defparam \D_iw[31] .power_up = "low";

cyclone10lp_lcell_comb \W_rf_wr_data[16]~11 (
	.dataa(\av_ld_byte2_data[0]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_16),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[16]~11_combout ),
	.cout());
defparam \W_rf_wr_data[16]~11 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[16]~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_rf_wr_data[15]~12 (
	.dataa(\av_ld_byte1_data[7]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_15),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[15]~12_combout ),
	.cout());
defparam \W_rf_wr_data[15]~12 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[15]~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_rf_wr_data[14]~13 (
	.dataa(\av_ld_byte1_data[6]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_14),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[14]~13_combout ),
	.cout());
defparam \W_rf_wr_data[14]~13 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[14]~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_rf_wr_data[13]~14 (
	.dataa(\av_ld_byte1_data[5]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_13),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[13]~14_combout ),
	.cout());
defparam \W_rf_wr_data[13]~14 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[13]~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_rf_wr_data[12]~15 (
	.dataa(\av_ld_byte1_data[4]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_12),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[12]~15_combout ),
	.cout());
defparam \W_rf_wr_data[12]~15 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[12]~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_rf_wr_data[11]~16 (
	.dataa(\av_ld_byte1_data[3]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_11),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[11]~16_combout ),
	.cout());
defparam \W_rf_wr_data[11]~16 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[11]~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_rf_wr_data[10]~17 (
	.dataa(\av_ld_byte1_data[2]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_10),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[10]~17_combout ),
	.cout());
defparam \W_rf_wr_data[10]~17 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[10]~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_rf_wr_data[9]~18 (
	.dataa(\av_ld_byte1_data[1]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_9),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[9]~18_combout ),
	.cout());
defparam \W_rf_wr_data[9]~18 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[9]~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_rf_wr_data[8]~19 (
	.dataa(\av_ld_byte1_data[0]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_8),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[8]~19_combout ),
	.cout());
defparam \W_rf_wr_data[8]~19 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[8]~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[1]~12 (
	.dataa(src0_valid),
	.datab(src0_valid1),
	.datac(av_readdata_pre_11),
	.datad(av_readdata_pre_1),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[1]~12_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[1]~12 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[1]~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[1]~13 (
	.dataa(read_latency_shift_reg_01),
	.datab(q_a_1),
	.datac(mem_74_01),
	.datad(mem_56_01),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[1]~13_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[1]~13 .lut_mask = 16'hEFFF;
defparam \av_ld_byte0_data_nxt[1]~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[1]~14 (
	.dataa(\av_ld_byte0_data_nxt[1]~12_combout ),
	.datab(\av_ld_byte0_data_nxt[1]~13_combout ),
	.datac(src0_valid3),
	.datad(av_readdata_pre_14),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[1]~14_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[1]~14 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[1]~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[1]~15 (
	.dataa(src0_valid5),
	.datab(src0_valid6),
	.datac(av_readdata_pre_12),
	.datad(av_readdata_pre_13),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[1]~15_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[1]~15 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[1]~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[1]~16 (
	.dataa(\av_ld_byte0_data_nxt[1]~15_combout ),
	.datab(src0_valid4),
	.datac(av_readdata_pre_15),
	.datad(gnd),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[1]~16_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[1]~16 .lut_mask = 16'hFEFE;
defparam \av_ld_byte0_data_nxt[1]~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[1]~17 (
	.dataa(\av_ld_byte1_data[1]~q ),
	.datab(\av_ld_byte0_data_nxt[1]~14_combout ),
	.datac(\av_ld_byte0_data_nxt[1]~16_combout ),
	.datad(\av_ld_rshift8~1_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[1]~17_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[1]~17 .lut_mask = 16'hFAFC;
defparam \av_ld_byte0_data_nxt[1]~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_control_rd_data[1]~4 (
	.dataa(\D_iw[8]~q ),
	.datab(\Equal135~0_combout ),
	.datac(\W_ipending_reg[1]~q ),
	.datad(\E_wrctl_status~0_combout ),
	.cin(gnd),
	.combout(\E_control_rd_data[1]~4_combout ),
	.cout());
defparam \E_control_rd_data[1]~4 .lut_mask = 16'hFFFE;
defparam \E_control_rd_data[1]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_control_rd_data[1]~5 (
	.dataa(\E_control_rd_data[1]~4_combout ),
	.datab(\Equal135~1_combout ),
	.datac(\W_ienable_reg[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\E_control_rd_data[1]~5_combout ),
	.cout());
defparam \E_control_rd_data[1]~5 .lut_mask = 16'hFEFE;
defparam \E_control_rd_data[1]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[2]~18 (
	.dataa(src0_valid),
	.datab(src0_valid1),
	.datac(av_readdata_pre_2),
	.datad(av_readdata_pre_27),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[2]~18_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[2]~18 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[2]~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[2]~19 (
	.dataa(read_latency_shift_reg_01),
	.datab(q_a_2),
	.datac(mem_74_01),
	.datad(mem_56_01),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[2]~19_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[2]~19 .lut_mask = 16'hEFFF;
defparam \av_ld_byte0_data_nxt[2]~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[2]~20 (
	.dataa(\av_ld_byte0_data_nxt[2]~18_combout ),
	.datab(\av_ld_byte0_data_nxt[2]~19_combout ),
	.datac(src0_valid4),
	.datad(av_readdata_pre_29),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[2]~20_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[2]~20 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[2]~20 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[2]~21 (
	.dataa(src0_valid5),
	.datab(src0_valid6),
	.datac(av_readdata_pre_210),
	.datad(av_readdata_pre_28),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[2]~21_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[2]~21 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[2]~21 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[2]~22 (
	.dataa(\av_ld_byte1_data[2]~q ),
	.datab(\av_ld_byte0_data_nxt[2]~20_combout ),
	.datac(\av_ld_byte0_data_nxt[2]~21_combout ),
	.datad(\av_ld_rshift8~1_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[2]~22_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[2]~22 .lut_mask = 16'hFAFC;
defparam \av_ld_byte0_data_nxt[2]~22 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[3]~23 (
	.dataa(src0_valid5),
	.datab(av_readdata_pre_33),
	.datac(src0_valid1),
	.datad(av_readdata_pre_31),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[3]~23_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[3]~23 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[3]~23 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[3]~24 (
	.dataa(src0_valid6),
	.datab(av_readdata_pre_32),
	.datac(src0_valid),
	.datad(av_readdata_pre_3),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[3]~24_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[3]~24 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[3]~24 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[3]~25 (
	.dataa(src0_valid2),
	.datab(q_a_3),
	.datac(\av_ld_byte0_data_nxt[3]~23_combout ),
	.datad(\av_ld_byte0_data_nxt[3]~24_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[3]~25_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[3]~25 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[3]~25 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[4]~26 (
	.dataa(src0_valid5),
	.datab(av_readdata_pre_4),
	.datac(src0_valid1),
	.datad(av_readdata_pre_42),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[4]~26_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[4]~26 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[4]~26 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[4]~27 (
	.dataa(src0_valid6),
	.datab(av_readdata_pre_41),
	.datac(src0_valid),
	.datad(av_readdata_pre_43),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[4]~27_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[4]~27 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[4]~27 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[4]~28 (
	.dataa(src0_valid2),
	.datab(q_a_4),
	.datac(\av_ld_byte0_data_nxt[4]~26_combout ),
	.datad(\av_ld_byte0_data_nxt[4]~27_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[4]~28_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[4]~28 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[4]~28 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[5]~29 (
	.dataa(src0_valid5),
	.datab(av_readdata_pre_5),
	.datac(src0_valid1),
	.datad(av_readdata_pre_52),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[5]~29_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[5]~29 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[5]~29 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[5]~30 (
	.dataa(src0_valid6),
	.datab(av_readdata_pre_51),
	.datac(src0_valid),
	.datad(av_readdata_pre_53),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[5]~30_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[5]~30 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[5]~30 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[5]~31 (
	.dataa(src0_valid2),
	.datab(q_a_5),
	.datac(\av_ld_byte0_data_nxt[5]~29_combout ),
	.datad(\av_ld_byte0_data_nxt[5]~30_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[5]~31_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[5]~31 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[5]~31 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[6]~32 (
	.dataa(src0_valid),
	.datab(src0_valid1),
	.datac(av_readdata_pre_6),
	.datad(av_readdata_pre_61),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[6]~32_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[6]~32 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[6]~32 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[6]~33 (
	.dataa(src0_valid2),
	.datab(src0_valid5),
	.datac(av_readdata_pre_62),
	.datad(q_a_6),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[6]~33_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[6]~33 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[6]~33 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[6]~34 (
	.dataa(\av_ld_byte0_data_nxt[6]~32_combout ),
	.datab(\av_ld_byte0_data_nxt[6]~33_combout ),
	.datac(src0_valid6),
	.datad(av_readdata_pre_63),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[6]~34_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[6]~34 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[6]~34 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[7]~35 (
	.dataa(src0_valid5),
	.datab(av_readdata_pre_72),
	.datac(src0_valid1),
	.datad(av_readdata_pre_7),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[7]~35_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[7]~35 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[7]~35 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[7]~36 (
	.dataa(src0_valid6),
	.datab(av_readdata_pre_73),
	.datac(src0_valid),
	.datad(av_readdata_pre_71),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[7]~36_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[7]~36 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[7]~36 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[7]~37 (
	.dataa(src0_valid2),
	.datab(q_a_7),
	.datac(\av_ld_byte0_data_nxt[7]~35_combout ),
	.datad(\av_ld_byte0_data_nxt[7]~36_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[7]~37_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[7]~37 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[7]~37 .sum_lutc_input = "datac";

dffeas R_ctrl_ld_signed(
	.clk(clk_clk),
	.d(\D_ctrl_ld_signed~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_ld_signed~q ),
	.prn(vcc));
defparam R_ctrl_ld_signed.is_wysiwyg = "true";
defparam R_ctrl_ld_signed.power_up = "low";

cyclone10lp_lcell_comb \av_fill_bit~0 (
	.dataa(\R_ctrl_ld_signed~q ),
	.datab(\av_ld_byte1_data[7]~q ),
	.datac(\av_ld_byte0_data[7]~q ),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\av_fill_bit~0_combout ),
	.cout());
defparam \av_fill_bit~0 .lut_mask = 16'hFAFC;
defparam \av_fill_bit~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte1_data_en~0 (
	.dataa(\D_iw[4]~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(\av_ld_aligning_data~q ),
	.datad(\D_ctrl_mem16~0_combout ),
	.cin(gnd),
	.combout(\av_ld_byte1_data_en~0_combout ),
	.cout());
defparam \av_ld_byte1_data_en~0 .lut_mask = 16'hEFFF;
defparam \av_ld_byte1_data_en~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[27]~73 (
	.dataa(read_latency_shift_reg_0),
	.datab(mem_74_0),
	.datac(mem_56_0),
	.datad(av_readdata_pre_271),
	.cin(gnd),
	.combout(\F_iw[27]~73_combout ),
	.cout());
defparam \F_iw[27]~73 .lut_mask = 16'hFFFE;
defparam \F_iw[27]~73 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[27]~74 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[27]~73_combout ),
	.datac(src1_valid2),
	.datad(q_a_27),
	.cin(gnd),
	.combout(\F_iw[27]~74_combout ),
	.cout());
defparam \F_iw[27]~74 .lut_mask = 16'hFFFE;
defparam \F_iw[27]~74 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[28]~75 (
	.dataa(read_latency_shift_reg_0),
	.datab(mem_74_0),
	.datac(mem_56_0),
	.datad(av_readdata_pre_281),
	.cin(gnd),
	.combout(\F_iw[28]~75_combout ),
	.cout());
defparam \F_iw[28]~75 .lut_mask = 16'hFFFE;
defparam \F_iw[28]~75 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[28]~76 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[28]~75_combout ),
	.datac(src1_valid2),
	.datad(q_a_28),
	.cin(gnd),
	.combout(\F_iw[28]~76_combout ),
	.cout());
defparam \F_iw[28]~76 .lut_mask = 16'hFFFE;
defparam \F_iw[28]~76 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[29]~77 (
	.dataa(read_latency_shift_reg_0),
	.datab(mem_74_0),
	.datac(mem_56_0),
	.datad(av_readdata_pre_291),
	.cin(gnd),
	.combout(\F_iw[29]~77_combout ),
	.cout());
defparam \F_iw[29]~77 .lut_mask = 16'hFFFE;
defparam \F_iw[29]~77 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[29]~78 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[29]~77_combout ),
	.datac(src1_valid2),
	.datad(q_a_29),
	.cin(gnd),
	.combout(\F_iw[29]~78_combout ),
	.cout());
defparam \F_iw[29]~78 .lut_mask = 16'hFFFE;
defparam \F_iw[29]~78 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[30]~79 (
	.dataa(read_latency_shift_reg_0),
	.datab(mem_74_0),
	.datac(mem_56_0),
	.datad(av_readdata_pre_30),
	.cin(gnd),
	.combout(\F_iw[30]~79_combout ),
	.cout());
defparam \F_iw[30]~79 .lut_mask = 16'hFFFE;
defparam \F_iw[30]~79 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[30]~80 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[30]~79_combout ),
	.datac(src1_valid2),
	.datad(q_a_30),
	.cin(gnd),
	.combout(\F_iw[30]~80_combout ),
	.cout());
defparam \F_iw[30]~80 .lut_mask = 16'hFFFE;
defparam \F_iw[30]~80 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[31]~81 (
	.dataa(read_latency_shift_reg_0),
	.datab(mem_74_0),
	.datac(mem_56_0),
	.datad(av_readdata_pre_311),
	.cin(gnd),
	.combout(\F_iw[31]~81_combout ),
	.cout());
defparam \F_iw[31]~81 .lut_mask = 16'hFFFE;
defparam \F_iw[31]~81 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[31]~82 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[31]~81_combout ),
	.datac(src1_valid2),
	.datad(q_a_31),
	.cin(gnd),
	.combout(\F_iw[31]~82_combout ),
	.cout());
defparam \F_iw[31]~82 .lut_mask = 16'hFFFE;
defparam \F_iw[31]~82 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[7] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[7]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[7] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[7] .power_up = "low";

cyclone10lp_lcell_comb \W_rf_wr_data[31]~20 (
	.dataa(\av_ld_byte3_data[7]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[31]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[31]~20_combout ),
	.cout());
defparam \W_rf_wr_data[31]~20 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[31]~20 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[6] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[6]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[6] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[6] .power_up = "low";

cyclone10lp_lcell_comb \W_rf_wr_data[30]~21 (
	.dataa(\av_ld_byte3_data[6]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[30]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[30]~21_combout ),
	.cout());
defparam \W_rf_wr_data[30]~21 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[30]~21 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[5] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[5]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[5] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[5] .power_up = "low";

cyclone10lp_lcell_comb \W_rf_wr_data[29]~22 (
	.dataa(\av_ld_byte3_data[5]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[29]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[29]~22_combout ),
	.cout());
defparam \W_rf_wr_data[29]~22 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[29]~22 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[4] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[4]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[4] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[4] .power_up = "low";

cyclone10lp_lcell_comb \W_rf_wr_data[28]~23 (
	.dataa(\av_ld_byte3_data[4]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[28]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[28]~23_combout ),
	.cout());
defparam \W_rf_wr_data[28]~23 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[28]~23 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[3] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[3]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[3] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[3] .power_up = "low";

cyclone10lp_lcell_comb \W_rf_wr_data[27]~24 (
	.dataa(\av_ld_byte3_data[3]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[27]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[27]~24_combout ),
	.cout());
defparam \W_rf_wr_data[27]~24 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[27]~24 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[2] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[2]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[2] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[2] .power_up = "low";

cyclone10lp_lcell_comb \W_rf_wr_data[26]~25 (
	.dataa(\av_ld_byte3_data[2]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[26]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[26]~25_combout ),
	.cout());
defparam \W_rf_wr_data[26]~25 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[26]~25 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[1] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[1]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[1] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[1] .power_up = "low";

cyclone10lp_lcell_comb \W_rf_wr_data[25]~26 (
	.dataa(\av_ld_byte3_data[1]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[25]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[25]~26_combout ),
	.cout());
defparam \W_rf_wr_data[25]~26 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[25]~26 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[0] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[0]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[0] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[0] .power_up = "low";

cyclone10lp_lcell_comb \W_rf_wr_data[24]~27 (
	.dataa(\av_ld_byte3_data[0]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[24]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[24]~27_combout ),
	.cout());
defparam \W_rf_wr_data[24]~27 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[24]~27 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_rf_wr_data[23]~28 (
	.dataa(\av_ld_byte2_data[7]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[23]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[23]~28_combout ),
	.cout());
defparam \W_rf_wr_data[23]~28 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[23]~28 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_rf_wr_data[22]~29 (
	.dataa(\av_ld_byte2_data[6]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[22]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[22]~29_combout ),
	.cout());
defparam \W_rf_wr_data[22]~29 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[22]~29 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_rf_wr_data[21]~30 (
	.dataa(\av_ld_byte2_data[5]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[21]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[21]~30_combout ),
	.cout());
defparam \W_rf_wr_data[21]~30 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[21]~30 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_rf_wr_data[20]~31 (
	.dataa(\av_ld_byte2_data[4]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[20]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[20]~31_combout ),
	.cout());
defparam \W_rf_wr_data[20]~31 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[20]~31 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_rf_wr_data[19]~32 (
	.dataa(\av_ld_byte2_data[3]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[19]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[19]~32_combout ),
	.cout());
defparam \W_rf_wr_data[19]~32 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[19]~32 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_rf_wr_data[18]~33 (
	.dataa(\av_ld_byte2_data[2]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[18]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[18]~33_combout ),
	.cout());
defparam \W_rf_wr_data[18]~33 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[18]~33 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_rf_wr_data[17]~34 (
	.dataa(\av_ld_byte2_data[1]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[17]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[17]~34_combout ),
	.cout());
defparam \W_rf_wr_data[17]~34 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[17]~34 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte3_data_nxt~0 (
	.dataa(src0_valid1),
	.datab(src0_valid2),
	.datac(q_a_31),
	.datad(av_readdata_pre_311),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~0_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~0 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte3_data_nxt~1 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~1_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~1 .lut_mask = 16'hAACC;
defparam \av_ld_byte3_data_nxt~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte3_data_nxt~2 (
	.dataa(src0_valid1),
	.datab(src0_valid2),
	.datac(q_a_30),
	.datad(av_readdata_pre_30),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~2_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~2 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte3_data_nxt~3 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~2_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~3_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~3 .lut_mask = 16'hAACC;
defparam \av_ld_byte3_data_nxt~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte3_data_nxt~4 (
	.dataa(src0_valid1),
	.datab(src0_valid2),
	.datac(q_a_29),
	.datad(av_readdata_pre_291),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~4_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~4 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte3_data_nxt~5 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~4_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~5_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~5 .lut_mask = 16'hAACC;
defparam \av_ld_byte3_data_nxt~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte3_data_nxt~6 (
	.dataa(src0_valid1),
	.datab(src0_valid2),
	.datac(q_a_28),
	.datad(av_readdata_pre_281),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~6_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~6 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte3_data_nxt~7 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~6_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~7_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~7 .lut_mask = 16'hAACC;
defparam \av_ld_byte3_data_nxt~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte3_data_nxt~8 (
	.dataa(src0_valid1),
	.datab(src0_valid2),
	.datac(q_a_27),
	.datad(av_readdata_pre_271),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~8_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~8 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte3_data_nxt~9 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~8_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~9_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~9 .lut_mask = 16'hAACC;
defparam \av_ld_byte3_data_nxt~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte3_data_nxt~10 (
	.dataa(src0_valid1),
	.datab(src0_valid2),
	.datac(q_a_26),
	.datad(av_readdata_pre_26),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~10_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~10 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte3_data_nxt~11 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~10_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~11_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~11 .lut_mask = 16'hAACC;
defparam \av_ld_byte3_data_nxt~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte3_data_nxt~12 (
	.dataa(src0_valid1),
	.datab(src0_valid2),
	.datac(q_a_25),
	.datad(av_readdata_pre_25),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~12_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~12 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte3_data_nxt~13 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~12_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~13_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~13 .lut_mask = 16'hAACC;
defparam \av_ld_byte3_data_nxt~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte3_data_nxt~14 (
	.dataa(src0_valid1),
	.datab(src0_valid2),
	.datac(q_a_24),
	.datad(av_readdata_pre_24),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~14_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~14 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte3_data_nxt~15 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~14_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~15_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~15 .lut_mask = 16'hAACC;
defparam \av_ld_byte3_data_nxt~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal0~23 (
	.dataa(\D_iw[4]~q ),
	.datab(\D_iw[5]~q ),
	.datac(\Equal0~7_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal0~23_combout ),
	.cout());
defparam \Equal0~23 .lut_mask = 16'hF7F7;
defparam \Equal0~23 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[0]~38 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(\av_ld_byte1_data[0]~q ),
	.datad(src_data_0),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[0]~38_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[0]~38 .lut_mask = 16'hFFF6;
defparam \av_ld_byte0_data_nxt[0]~38 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_dst_regnum[1]~11 (
	.dataa(\D_iw[4]~q ),
	.datab(\D_iw[5]~q ),
	.datac(\Equal0~7_combout ),
	.datad(\D_dst_regnum[1]~3_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[1]~11_combout ),
	.cout());
defparam \D_dst_regnum[1]~11 .lut_mask = 16'hFFF7;
defparam \D_dst_regnum[1]~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[3]~39 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(\av_ld_byte1_data[3]~q ),
	.datad(\av_ld_byte0_data_nxt[3]~25_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[3]~39_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[3]~39 .lut_mask = 16'hFFF6;
defparam \av_ld_byte0_data_nxt[3]~39 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[4]~40 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(\av_ld_byte1_data[4]~q ),
	.datad(\av_ld_byte0_data_nxt[4]~28_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[4]~40_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[4]~40 .lut_mask = 16'hFFF6;
defparam \av_ld_byte0_data_nxt[4]~40 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[5]~41 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(\av_ld_byte1_data[5]~q ),
	.datad(\av_ld_byte0_data_nxt[5]~31_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[5]~41_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[5]~41 .lut_mask = 16'hFFF6;
defparam \av_ld_byte0_data_nxt[5]~41 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[6]~42 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(\av_ld_byte1_data[6]~q ),
	.datad(\av_ld_byte0_data_nxt[6]~34_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[6]~42_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[6]~42 .lut_mask = 16'hFFF6;
defparam \av_ld_byte0_data_nxt[6]~42 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_byte0_data_nxt[7]~43 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(\av_ld_byte1_data[7]~q ),
	.datad(\av_ld_byte0_data_nxt[7]~37_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[7]~43_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[7]~43 .lut_mask = 16'hFFF6;
defparam \av_ld_byte0_data_nxt[7]~43 .sum_lutc_input = "datac";

dffeas \W_alu_result[7] (
	.clk(clk_clk),
	.d(\W_alu_result[7]~9_combout ),
	.asdata(\E_shift_rot_result[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_7),
	.prn(vcc));
defparam \W_alu_result[7] .is_wysiwyg = "true";
defparam \W_alu_result[7] .power_up = "low";

dffeas \W_alu_result[16] (
	.clk(clk_clk),
	.d(\W_alu_result[16]~0_combout ),
	.asdata(\E_shift_rot_result[16]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_16),
	.prn(vcc));
defparam \W_alu_result[16] .is_wysiwyg = "true";
defparam \W_alu_result[16] .power_up = "low";

dffeas \W_alu_result[15] (
	.clk(clk_clk),
	.d(\W_alu_result[15]~1_combout ),
	.asdata(\E_shift_rot_result[15]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_15),
	.prn(vcc));
defparam \W_alu_result[15] .is_wysiwyg = "true";
defparam \W_alu_result[15] .power_up = "low";

dffeas \W_alu_result[14] (
	.clk(clk_clk),
	.d(\W_alu_result[14]~2_combout ),
	.asdata(\E_shift_rot_result[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_14),
	.prn(vcc));
defparam \W_alu_result[14] .is_wysiwyg = "true";
defparam \W_alu_result[14] .power_up = "low";

dffeas \W_alu_result[13] (
	.clk(clk_clk),
	.d(\W_alu_result[13]~3_combout ),
	.asdata(\E_shift_rot_result[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_13),
	.prn(vcc));
defparam \W_alu_result[13] .is_wysiwyg = "true";
defparam \W_alu_result[13] .power_up = "low";

dffeas \W_alu_result[12] (
	.clk(clk_clk),
	.d(\W_alu_result[12]~4_combout ),
	.asdata(\E_shift_rot_result[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_12),
	.prn(vcc));
defparam \W_alu_result[12] .is_wysiwyg = "true";
defparam \W_alu_result[12] .power_up = "low";

dffeas \W_alu_result[11] (
	.clk(clk_clk),
	.d(\W_alu_result[11]~5_combout ),
	.asdata(\E_shift_rot_result[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_11),
	.prn(vcc));
defparam \W_alu_result[11] .is_wysiwyg = "true";
defparam \W_alu_result[11] .power_up = "low";

dffeas \W_alu_result[10] (
	.clk(clk_clk),
	.d(\W_alu_result[10]~6_combout ),
	.asdata(\E_shift_rot_result[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_10),
	.prn(vcc));
defparam \W_alu_result[10] .is_wysiwyg = "true";
defparam \W_alu_result[10] .power_up = "low";

dffeas \W_alu_result[9] (
	.clk(clk_clk),
	.d(\W_alu_result[9]~7_combout ),
	.asdata(\E_shift_rot_result[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_9),
	.prn(vcc));
defparam \W_alu_result[9] .is_wysiwyg = "true";
defparam \W_alu_result[9] .power_up = "low";

dffeas \W_alu_result[8] (
	.clk(clk_clk),
	.d(\W_alu_result[8]~8_combout ),
	.asdata(\E_shift_rot_result[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_8),
	.prn(vcc));
defparam \W_alu_result[8] .is_wysiwyg = "true";
defparam \W_alu_result[8] .power_up = "low";

dffeas \W_alu_result[4] (
	.clk(clk_clk),
	.d(\W_alu_result[4]~12_combout ),
	.asdata(\E_shift_rot_result[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_4),
	.prn(vcc));
defparam \W_alu_result[4] .is_wysiwyg = "true";
defparam \W_alu_result[4] .power_up = "low";

dffeas \W_alu_result[5] (
	.clk(clk_clk),
	.d(\W_alu_result[5]~11_combout ),
	.asdata(\E_shift_rot_result[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_5),
	.prn(vcc));
defparam \W_alu_result[5] .is_wysiwyg = "true";
defparam \W_alu_result[5] .power_up = "low";

dffeas \W_alu_result[6] (
	.clk(clk_clk),
	.d(\W_alu_result[6]~10_combout ),
	.asdata(\E_shift_rot_result[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_6),
	.prn(vcc));
defparam \W_alu_result[6] .is_wysiwyg = "true";
defparam \W_alu_result[6] .power_up = "low";

dffeas \W_alu_result[2] (
	.clk(clk_clk),
	.d(\W_alu_result[2]~13_combout ),
	.asdata(\E_shift_rot_result[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_2),
	.prn(vcc));
defparam \W_alu_result[2] .is_wysiwyg = "true";
defparam \W_alu_result[2] .power_up = "low";

dffeas \W_alu_result[3] (
	.clk(clk_clk),
	.d(\W_alu_result[3]~14_combout ),
	.asdata(\E_shift_rot_result[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_3),
	.prn(vcc));
defparam \W_alu_result[3] .is_wysiwyg = "true";
defparam \W_alu_result[3] .power_up = "low";

dffeas \d_writedata[24] (
	.clk(clk_clk),
	.d(\d_writedata[24]~0_combout ),
	.asdata(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_24),
	.prn(vcc));
defparam \d_writedata[24] .is_wysiwyg = "true";
defparam \d_writedata[24] .power_up = "low";

dffeas \d_writedata[25] (
	.clk(clk_clk),
	.d(\d_writedata[25]~1_combout ),
	.asdata(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_25),
	.prn(vcc));
defparam \d_writedata[25] .is_wysiwyg = "true";
defparam \d_writedata[25] .power_up = "low";

dffeas \d_writedata[26] (
	.clk(clk_clk),
	.d(\d_writedata[26]~2_combout ),
	.asdata(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_26),
	.prn(vcc));
defparam \d_writedata[26] .is_wysiwyg = "true";
defparam \d_writedata[26] .power_up = "low";

dffeas \d_writedata[27] (
	.clk(clk_clk),
	.d(\d_writedata[27]~3_combout ),
	.asdata(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_27),
	.prn(vcc));
defparam \d_writedata[27] .is_wysiwyg = "true";
defparam \d_writedata[27] .power_up = "low";

dffeas \d_writedata[28] (
	.clk(clk_clk),
	.d(\d_writedata[28]~4_combout ),
	.asdata(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_28),
	.prn(vcc));
defparam \d_writedata[28] .is_wysiwyg = "true";
defparam \d_writedata[28] .power_up = "low";

dffeas \d_writedata[29] (
	.clk(clk_clk),
	.d(\d_writedata[29]~5_combout ),
	.asdata(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_29),
	.prn(vcc));
defparam \d_writedata[29] .is_wysiwyg = "true";
defparam \d_writedata[29] .power_up = "low";

dffeas \d_writedata[30] (
	.clk(clk_clk),
	.d(\d_writedata[30]~6_combout ),
	.asdata(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_30),
	.prn(vcc));
defparam \d_writedata[30] .is_wysiwyg = "true";
defparam \d_writedata[30] .power_up = "low";

dffeas \d_writedata[31] (
	.clk(clk_clk),
	.d(\d_writedata[31]~7_combout ),
	.asdata(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_31),
	.prn(vcc));
defparam \d_writedata[31] .is_wysiwyg = "true";
defparam \d_writedata[31] .power_up = "low";

dffeas \d_writedata[0] (
	.clk(clk_clk),
	.d(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_0),
	.prn(vcc));
defparam \d_writedata[0] .is_wysiwyg = "true";
defparam \d_writedata[0] .power_up = "low";

dffeas d_write(
	.clk(clk_clk),
	.d(\E_st_stall~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_write1),
	.prn(vcc));
defparam d_write.is_wysiwyg = "true";
defparam d_write.power_up = "low";

dffeas i_read(
	.clk(clk_clk),
	.d(\i_read_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(i_read1),
	.prn(vcc));
defparam i_read.is_wysiwyg = "true";
defparam i_read.power_up = "low";

dffeas \F_pc[5] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[5]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_5),
	.prn(vcc));
defparam \F_pc[5] .is_wysiwyg = "true";
defparam \F_pc[5] .power_up = "low";

dffeas \F_pc[14] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[14]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_14),
	.prn(vcc));
defparam \F_pc[14] .is_wysiwyg = "true";
defparam \F_pc[14] .power_up = "low";

dffeas \F_pc[13] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[13]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_13),
	.prn(vcc));
defparam \F_pc[13] .is_wysiwyg = "true";
defparam \F_pc[13] .power_up = "low";

dffeas \F_pc[12] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[12]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_12),
	.prn(vcc));
defparam \F_pc[12] .is_wysiwyg = "true";
defparam \F_pc[12] .power_up = "low";

dffeas \F_pc[11] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[11]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_11),
	.prn(vcc));
defparam \F_pc[11] .is_wysiwyg = "true";
defparam \F_pc[11] .power_up = "low";

dffeas \F_pc[10] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[10]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_10),
	.prn(vcc));
defparam \F_pc[10] .is_wysiwyg = "true";
defparam \F_pc[10] .power_up = "low";

dffeas \F_pc[9] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[9]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_9),
	.prn(vcc));
defparam \F_pc[9] .is_wysiwyg = "true";
defparam \F_pc[9] .power_up = "low";

dffeas \F_pc[8] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[8]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_8),
	.prn(vcc));
defparam \F_pc[8] .is_wysiwyg = "true";
defparam \F_pc[8] .power_up = "low";

dffeas \F_pc[7] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[7]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_7),
	.prn(vcc));
defparam \F_pc[7] .is_wysiwyg = "true";
defparam \F_pc[7] .power_up = "low";

dffeas \F_pc[6] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[6]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_6),
	.prn(vcc));
defparam \F_pc[6] .is_wysiwyg = "true";
defparam \F_pc[6] .power_up = "low";

dffeas \F_pc[2] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[2]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_2),
	.prn(vcc));
defparam \F_pc[2] .is_wysiwyg = "true";
defparam \F_pc[2] .power_up = "low";

dffeas \F_pc[3] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[3]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_3),
	.prn(vcc));
defparam \F_pc[3] .is_wysiwyg = "true";
defparam \F_pc[3] .power_up = "low";

dffeas \F_pc[4] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[4]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_4),
	.prn(vcc));
defparam \F_pc[4] .is_wysiwyg = "true";
defparam \F_pc[4] .power_up = "low";

dffeas d_read(
	.clk(clk_clk),
	.d(\d_read_nxt~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_read1),
	.prn(vcc));
defparam d_read.is_wysiwyg = "true";
defparam d_read.power_up = "low";

dffeas \F_pc[1] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[1]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_1),
	.prn(vcc));
defparam \F_pc[1] .is_wysiwyg = "true";
defparam \F_pc[1] .power_up = "low";

dffeas \F_pc[0] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[0]~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_0),
	.prn(vcc));
defparam \F_pc[0] .is_wysiwyg = "true";
defparam \F_pc[0] .power_up = "low";

dffeas \d_writedata[1] (
	.clk(clk_clk),
	.d(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_1),
	.prn(vcc));
defparam \d_writedata[1] .is_wysiwyg = "true";
defparam \d_writedata[1] .power_up = "low";

dffeas \d_writedata[2] (
	.clk(clk_clk),
	.d(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_2),
	.prn(vcc));
defparam \d_writedata[2] .is_wysiwyg = "true";
defparam \d_writedata[2] .power_up = "low";

dffeas \d_writedata[3] (
	.clk(clk_clk),
	.d(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_3),
	.prn(vcc));
defparam \d_writedata[3] .is_wysiwyg = "true";
defparam \d_writedata[3] .power_up = "low";

dffeas \d_writedata[4] (
	.clk(clk_clk),
	.d(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_4),
	.prn(vcc));
defparam \d_writedata[4] .is_wysiwyg = "true";
defparam \d_writedata[4] .power_up = "low";

dffeas \d_writedata[5] (
	.clk(clk_clk),
	.d(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_5),
	.prn(vcc));
defparam \d_writedata[5] .is_wysiwyg = "true";
defparam \d_writedata[5] .power_up = "low";

dffeas \d_writedata[6] (
	.clk(clk_clk),
	.d(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_6),
	.prn(vcc));
defparam \d_writedata[6] .is_wysiwyg = "true";
defparam \d_writedata[6] .power_up = "low";

dffeas \d_writedata[7] (
	.clk(clk_clk),
	.d(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_7),
	.prn(vcc));
defparam \d_writedata[7] .is_wysiwyg = "true";
defparam \d_writedata[7] .power_up = "low";

dffeas \d_writedata[9] (
	.clk(clk_clk),
	.d(\E_st_data[9]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_9),
	.prn(vcc));
defparam \d_writedata[9] .is_wysiwyg = "true";
defparam \d_writedata[9] .power_up = "low";

dffeas hbreak_enabled(
	.clk(clk_clk),
	.d(\hbreak_enabled~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\E_valid_from_R~q ),
	.q(hbreak_enabled1),
	.prn(vcc));
defparam hbreak_enabled.is_wysiwyg = "true";
defparam hbreak_enabled.power_up = "low";

dffeas \d_byteenable[0] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_0),
	.prn(vcc));
defparam \d_byteenable[0] .is_wysiwyg = "true";
defparam \d_byteenable[0] .power_up = "low";

dffeas \d_writedata[22] (
	.clk(clk_clk),
	.d(\E_st_data[22]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_22),
	.prn(vcc));
defparam \d_writedata[22] .is_wysiwyg = "true";
defparam \d_writedata[22] .power_up = "low";

dffeas \d_byteenable[2] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[2]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_2),
	.prn(vcc));
defparam \d_byteenable[2] .is_wysiwyg = "true";
defparam \d_byteenable[2] .power_up = "low";

dffeas \d_writedata[23] (
	.clk(clk_clk),
	.d(\E_st_data[23]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_23),
	.prn(vcc));
defparam \d_writedata[23] .is_wysiwyg = "true";
defparam \d_writedata[23] .power_up = "low";

dffeas \d_byteenable[3] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[3]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_3),
	.prn(vcc));
defparam \d_byteenable[3] .is_wysiwyg = "true";
defparam \d_byteenable[3] .power_up = "low";

dffeas \d_writedata[14] (
	.clk(clk_clk),
	.d(\E_st_data[14]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_14),
	.prn(vcc));
defparam \d_writedata[14] .is_wysiwyg = "true";
defparam \d_writedata[14] .power_up = "low";

dffeas \d_byteenable[1] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[1]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_1),
	.prn(vcc));
defparam \d_byteenable[1] .is_wysiwyg = "true";
defparam \d_byteenable[1] .power_up = "low";

dffeas \d_writedata[15] (
	.clk(clk_clk),
	.d(\E_st_data[15]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_15),
	.prn(vcc));
defparam \d_writedata[15] .is_wysiwyg = "true";
defparam \d_writedata[15] .power_up = "low";

dffeas \d_writedata[11] (
	.clk(clk_clk),
	.d(\E_st_data[11]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_11),
	.prn(vcc));
defparam \d_writedata[11] .is_wysiwyg = "true";
defparam \d_writedata[11] .power_up = "low";

dffeas \d_writedata[13] (
	.clk(clk_clk),
	.d(\E_st_data[13]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_13),
	.prn(vcc));
defparam \d_writedata[13] .is_wysiwyg = "true";
defparam \d_writedata[13] .power_up = "low";

dffeas \d_writedata[16] (
	.clk(clk_clk),
	.d(\E_st_data[16]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_16),
	.prn(vcc));
defparam \d_writedata[16] .is_wysiwyg = "true";
defparam \d_writedata[16] .power_up = "low";

dffeas \d_writedata[12] (
	.clk(clk_clk),
	.d(\E_st_data[12]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_12),
	.prn(vcc));
defparam \d_writedata[12] .is_wysiwyg = "true";
defparam \d_writedata[12] .power_up = "low";

dffeas \d_writedata[10] (
	.clk(clk_clk),
	.d(\E_st_data[10]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_10),
	.prn(vcc));
defparam \d_writedata[10] .is_wysiwyg = "true";
defparam \d_writedata[10] .power_up = "low";

dffeas \d_writedata[8] (
	.clk(clk_clk),
	.d(\E_st_data[8]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_8),
	.prn(vcc));
defparam \d_writedata[8] .is_wysiwyg = "true";
defparam \d_writedata[8] .power_up = "low";

dffeas \d_writedata[21] (
	.clk(clk_clk),
	.d(\E_st_data[21]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_21),
	.prn(vcc));
defparam \d_writedata[21] .is_wysiwyg = "true";
defparam \d_writedata[21] .power_up = "low";

dffeas \d_writedata[20] (
	.clk(clk_clk),
	.d(\E_st_data[20]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_20),
	.prn(vcc));
defparam \d_writedata[20] .is_wysiwyg = "true";
defparam \d_writedata[20] .power_up = "low";

dffeas \d_writedata[19] (
	.clk(clk_clk),
	.d(\E_st_data[19]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_19),
	.prn(vcc));
defparam \d_writedata[19] .is_wysiwyg = "true";
defparam \d_writedata[19] .power_up = "low";

dffeas \d_writedata[18] (
	.clk(clk_clk),
	.d(\E_st_data[18]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_18),
	.prn(vcc));
defparam \d_writedata[18] .is_wysiwyg = "true";
defparam \d_writedata[18] .power_up = "low";

dffeas \d_writedata[17] (
	.clk(clk_clk),
	.d(\E_st_data[17]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_17),
	.prn(vcc));
defparam \d_writedata[17] .is_wysiwyg = "true";
defparam \d_writedata[17] .power_up = "low";

cyclone10lp_lcell_comb \F_valid~0 (
	.dataa(WideOr13),
	.datab(WideOr14),
	.datac(gnd),
	.datad(i_read1),
	.cin(gnd),
	.combout(\F_valid~0_combout ),
	.cout());
defparam \F_valid~0 .lut_mask = 16'hEEFF;
defparam \F_valid~0 .sum_lutc_input = "datac";

dffeas D_valid(
	.clk(clk_clk),
	.d(\F_valid~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\D_valid~q ),
	.prn(vcc));
defparam D_valid.is_wysiwyg = "true";
defparam D_valid.power_up = "low";

dffeas R_valid(
	.clk(clk_clk),
	.d(\D_valid~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_valid~q ),
	.prn(vcc));
defparam R_valid.is_wysiwyg = "true";
defparam R_valid.power_up = "low";

dffeas E_new_inst(
	.clk(clk_clk),
	.d(\R_valid~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_new_inst~q ),
	.prn(vcc));
defparam E_new_inst.is_wysiwyg = "true";
defparam E_new_inst.power_up = "low";

cyclone10lp_lcell_comb \F_iw[0]~14 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(src_data_01),
	.datac(src_data_02),
	.datad(src_data_03),
	.cin(gnd),
	.combout(\F_iw[0]~14_combout ),
	.cout());
defparam \F_iw[0]~14 .lut_mask = 16'hFFFE;
defparam \F_iw[0]~14 .sum_lutc_input = "datac";

dffeas \D_iw[0] (
	.clk(clk_clk),
	.d(\F_iw[0]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[0]~q ),
	.prn(vcc));
defparam \D_iw[0] .is_wysiwyg = "true";
defparam \D_iw[0] .power_up = "low";

cyclone10lp_lcell_comb \F_iw[4]~20 (
	.dataa(read_latency_shift_reg_02),
	.datab(mem_74_02),
	.datac(mem_56_02),
	.datad(av_readdata_pre_4),
	.cin(gnd),
	.combout(\F_iw[4]~20_combout ),
	.cout());
defparam \F_iw[4]~20 .lut_mask = 16'hFFFE;
defparam \F_iw[4]~20 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[4]~21 (
	.dataa(src1_valid4),
	.datab(av_readdata_pre_41),
	.datac(src1_valid1),
	.datad(av_readdata_pre_42),
	.cin(gnd),
	.combout(\F_iw[4]~21_combout ),
	.cout());
defparam \F_iw[4]~21 .lut_mask = 16'hFFFE;
defparam \F_iw[4]~21 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[4]~22 (
	.dataa(src1_valid2),
	.datab(q_a_4),
	.datac(\F_iw[4]~20_combout ),
	.datad(\F_iw[4]~21_combout ),
	.cin(gnd),
	.combout(\F_iw[4]~22_combout ),
	.cout());
defparam \F_iw[4]~22 .lut_mask = 16'hFFFE;
defparam \F_iw[4]~22 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[4]~23 (
	.dataa(\F_iw[4]~22_combout ),
	.datab(src1_valid),
	.datac(av_readdata_pre_43),
	.datad(\D_iw[26]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[4]~23_combout ),
	.cout());
defparam \F_iw[4]~23 .lut_mask = 16'hFEFF;
defparam \F_iw[4]~23 .sum_lutc_input = "datac";

dffeas \D_iw[4] (
	.clk(clk_clk),
	.d(\F_iw[4]~23_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[4]~q ),
	.prn(vcc));
defparam \D_iw[4] .is_wysiwyg = "true";
defparam \D_iw[4] .power_up = "low";

cyclone10lp_lcell_comb \F_iw[3]~24 (
	.dataa(src1_valid1),
	.datab(src1_valid2),
	.datac(q_a_3),
	.datad(av_readdata_pre_31),
	.cin(gnd),
	.combout(\F_iw[3]~24_combout ),
	.cout());
defparam \F_iw[3]~24 .lut_mask = 16'hFFFE;
defparam \F_iw[3]~24 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[3]~25 (
	.dataa(src1_valid3),
	.datab(src1_valid4),
	.datac(av_readdata_pre_32),
	.datad(av_readdata_pre_33),
	.cin(gnd),
	.combout(\F_iw[3]~25_combout ),
	.cout());
defparam \F_iw[3]~25 .lut_mask = 16'hFFFE;
defparam \F_iw[3]~25 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[3]~26 (
	.dataa(src_payload2),
	.datab(\F_iw[3]~24_combout ),
	.datac(\F_iw[3]~25_combout ),
	.datad(\D_iw[26]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[3]~26_combout ),
	.cout());
defparam \F_iw[3]~26 .lut_mask = 16'hFEFF;
defparam \F_iw[3]~26 .sum_lutc_input = "datac";

dffeas \D_iw[3] (
	.clk(clk_clk),
	.d(\F_iw[3]~26_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[3]~q ),
	.prn(vcc));
defparam \D_iw[3] .is_wysiwyg = "true";
defparam \D_iw[3] .power_up = "low";

cyclone10lp_lcell_comb \D_ctrl_st~0 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[4]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_st~0_combout ),
	.cout());
defparam \D_ctrl_st~0 .lut_mask = 16'hBFFF;
defparam \D_ctrl_st~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[2]~27 (
	.dataa(src1_valid),
	.datab(src1_valid1),
	.datac(av_readdata_pre_2),
	.datad(av_readdata_pre_27),
	.cin(gnd),
	.combout(\F_iw[2]~27_combout ),
	.cout());
defparam \F_iw[2]~27 .lut_mask = 16'hFFFE;
defparam \F_iw[2]~27 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[2]~28 (
	.dataa(src1_valid2),
	.datab(src1_valid3),
	.datac(av_readdata_pre_28),
	.datad(q_a_2),
	.cin(gnd),
	.combout(\F_iw[2]~28_combout ),
	.cout());
defparam \F_iw[2]~28 .lut_mask = 16'hFFFE;
defparam \F_iw[2]~28 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[2]~29 (
	.dataa(src1_valid4),
	.datab(src_payload),
	.datac(av_readdata_pre_29),
	.datad(av_readdata_pre_210),
	.cin(gnd),
	.combout(\F_iw[2]~29_combout ),
	.cout());
defparam \F_iw[2]~29 .lut_mask = 16'hFFFE;
defparam \F_iw[2]~29 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[2]~30 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[2]~27_combout ),
	.datac(\F_iw[2]~28_combout ),
	.datad(\F_iw[2]~29_combout ),
	.cin(gnd),
	.combout(\F_iw[2]~30_combout ),
	.cout());
defparam \F_iw[2]~30 .lut_mask = 16'hFFFE;
defparam \F_iw[2]~30 .sum_lutc_input = "datac";

dffeas \D_iw[2] (
	.clk(clk_clk),
	.d(\F_iw[2]~30_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[2]~q ),
	.prn(vcc));
defparam \D_iw[2] .is_wysiwyg = "true";
defparam \D_iw[2] .power_up = "low";

dffeas R_ctrl_st(
	.clk(clk_clk),
	.d(\D_ctrl_st~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!\D_iw[2]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_st~q ),
	.prn(vcc));
defparam R_ctrl_st.is_wysiwyg = "true";
defparam R_ctrl_st.power_up = "low";

cyclone10lp_lcell_comb E_st_stall(
	.dataa(d_write1),
	.datab(\E_new_inst~q ),
	.datac(\R_ctrl_st~q ),
	.datad(av_waitrequest),
	.cin(gnd),
	.combout(\E_st_stall~combout ),
	.cout());
defparam E_st_stall.lut_mask = 16'hFFFE;
defparam E_st_stall.sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[5]~31 (
	.dataa(read_latency_shift_reg_02),
	.datab(mem_74_02),
	.datac(mem_56_02),
	.datad(av_readdata_pre_5),
	.cin(gnd),
	.combout(\F_iw[5]~31_combout ),
	.cout());
defparam \F_iw[5]~31 .lut_mask = 16'hFFFE;
defparam \F_iw[5]~31 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[5]~32 (
	.dataa(src1_valid4),
	.datab(av_readdata_pre_51),
	.datac(src1_valid1),
	.datad(av_readdata_pre_52),
	.cin(gnd),
	.combout(\F_iw[5]~32_combout ),
	.cout());
defparam \F_iw[5]~32 .lut_mask = 16'hFFFE;
defparam \F_iw[5]~32 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[5]~33 (
	.dataa(src1_valid2),
	.datab(q_a_5),
	.datac(\F_iw[5]~31_combout ),
	.datad(\F_iw[5]~32_combout ),
	.cin(gnd),
	.combout(\F_iw[5]~33_combout ),
	.cout());
defparam \F_iw[5]~33 .lut_mask = 16'hFFFE;
defparam \F_iw[5]~33 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[5]~34 (
	.dataa(\F_iw[5]~33_combout ),
	.datab(src1_valid),
	.datac(av_readdata_pre_53),
	.datad(\D_iw[26]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[5]~34_combout ),
	.cout());
defparam \F_iw[5]~34 .lut_mask = 16'hFEFF;
defparam \F_iw[5]~34 .sum_lutc_input = "datac";

dffeas \D_iw[5] (
	.clk(clk_clk),
	.d(\F_iw[5]~34_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[5]~q ),
	.prn(vcc));
defparam \D_iw[5] .is_wysiwyg = "true";
defparam \D_iw[5] .power_up = "low";

cyclone10lp_lcell_comb \Equal0~9 (
	.dataa(\D_iw[4]~q ),
	.datab(\Equal0~4_combout ),
	.datac(\D_iw[5]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal0~9_combout ),
	.cout());
defparam \Equal0~9 .lut_mask = 16'hFEFE;
defparam \Equal0~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_valid~0 (
	.dataa(\E_valid_from_R~q ),
	.datab(gnd),
	.datac(\E_st_stall~combout ),
	.datad(\E_stall~4_combout ),
	.cin(gnd),
	.combout(\W_valid~0_combout ),
	.cout());
defparam \W_valid~0 .lut_mask = 16'hAFFF;
defparam \W_valid~0 .sum_lutc_input = "datac";

dffeas W_valid(
	.clk(clk_clk),
	.d(\W_valid~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_valid~q ),
	.prn(vcc));
defparam W_valid.is_wysiwyg = "true";
defparam W_valid.power_up = "low";

cyclone10lp_lcell_comb \hbreak_pending_nxt~0 (
	.dataa(\hbreak_pending~q ),
	.datab(\hbreak_req~0_combout ),
	.datac(gnd),
	.datad(hbreak_enabled1),
	.cin(gnd),
	.combout(\hbreak_pending_nxt~0_combout ),
	.cout());
defparam \hbreak_pending_nxt~0 .lut_mask = 16'hEEFF;
defparam \hbreak_pending_nxt~0 .sum_lutc_input = "datac";

dffeas hbreak_pending(
	.clk(clk_clk),
	.d(\hbreak_pending_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\hbreak_pending~q ),
	.prn(vcc));
defparam hbreak_pending.is_wysiwyg = "true";
defparam hbreak_pending.power_up = "low";

cyclone10lp_lcell_comb \wait_for_one_post_bret_inst~0 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_oci|the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_single_step_mode~q ),
	.datab(hbreak_enabled1),
	.datac(\wait_for_one_post_bret_inst~q ),
	.datad(\F_valid~0_combout ),
	.cin(gnd),
	.combout(\wait_for_one_post_bret_inst~0_combout ),
	.cout());
defparam \wait_for_one_post_bret_inst~0 .lut_mask = 16'hFEFF;
defparam \wait_for_one_post_bret_inst~0 .sum_lutc_input = "datac";

dffeas wait_for_one_post_bret_inst(
	.clk(clk_clk),
	.d(\wait_for_one_post_bret_inst~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wait_for_one_post_bret_inst~q ),
	.prn(vcc));
defparam wait_for_one_post_bret_inst.is_wysiwyg = "true";
defparam wait_for_one_post_bret_inst.power_up = "low";

cyclone10lp_lcell_comb \hbreak_req~0 (
	.dataa(\W_valid~q ),
	.datab(\hbreak_pending~q ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_oci|the_processor_nios2_gen2_0_cpu_nios2_oci_debug|jtag_break~q ),
	.datad(\wait_for_one_post_bret_inst~q ),
	.cin(gnd),
	.combout(\hbreak_req~0_combout ),
	.cout());
defparam \hbreak_req~0 .lut_mask = 16'hFEFF;
defparam \hbreak_req~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[14]~35 (
	.dataa(src1_valid1),
	.datab(src1_valid2),
	.datac(q_a_14),
	.datad(av_readdata_pre_141),
	.cin(gnd),
	.combout(\F_iw[14]~35_combout ),
	.cout());
defparam \F_iw[14]~35 .lut_mask = 16'hFFFE;
defparam \F_iw[14]~35 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[14]~36 (
	.dataa(\F_iw[14]~35_combout ),
	.datab(src1_valid),
	.datac(av_readdata_pre_142),
	.datad(gnd),
	.cin(gnd),
	.combout(\F_iw[14]~36_combout ),
	.cout());
defparam \F_iw[14]~36 .lut_mask = 16'hFEFE;
defparam \F_iw[14]~36 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[14]~83 (
	.dataa(\D_iw[26]~0_combout ),
	.datab(hbreak_enabled1),
	.datac(\hbreak_req~0_combout ),
	.datad(\F_iw[14]~36_combout ),
	.cin(gnd),
	.combout(\F_iw[14]~83_combout ),
	.cout());
defparam \F_iw[14]~83 .lut_mask = 16'hFFDF;
defparam \F_iw[14]~83 .sum_lutc_input = "datac";

dffeas \D_iw[14] (
	.clk(clk_clk),
	.d(\F_iw[14]~83_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[14]~q ),
	.prn(vcc));
defparam \D_iw[14] .is_wysiwyg = "true";
defparam \D_iw[14] .power_up = "low";

cyclone10lp_lcell_comb \F_iw[15]~37 (
	.dataa(src1_valid1),
	.datab(src1_valid2),
	.datac(q_a_15),
	.datad(av_readdata_pre_151),
	.cin(gnd),
	.combout(\F_iw[15]~37_combout ),
	.cout());
defparam \F_iw[15]~37 .lut_mask = 16'hFFFE;
defparam \F_iw[15]~37 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[15]~38 (
	.dataa(\F_iw[15]~37_combout ),
	.datab(src1_valid),
	.datac(av_readdata_pre_152),
	.datad(\D_iw[26]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[15]~38_combout ),
	.cout());
defparam \F_iw[15]~38 .lut_mask = 16'hFEFF;
defparam \F_iw[15]~38 .sum_lutc_input = "datac";

dffeas \D_iw[15] (
	.clk(clk_clk),
	.d(\F_iw[15]~38_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[15]~q ),
	.prn(vcc));
defparam \D_iw[15] .is_wysiwyg = "true";
defparam \D_iw[15] .power_up = "low";

cyclone10lp_lcell_comb \D_op_opx_rsv63~0 (
	.dataa(\D_iw[14]~q ),
	.datab(\D_iw[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_op_opx_rsv63~0_combout ),
	.cout());
defparam \D_op_opx_rsv63~0 .lut_mask = 16'hEEEE;
defparam \D_op_opx_rsv63~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[11]~39 (
	.dataa(src_payload3),
	.datab(src1_valid1),
	.datac(av_readdata_pre_111),
	.datad(\D_iw[26]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[11]~39_combout ),
	.cout());
defparam \F_iw[11]~39 .lut_mask = 16'hFEFF;
defparam \F_iw[11]~39 .sum_lutc_input = "datac";

dffeas \D_iw[11] (
	.clk(clk_clk),
	.d(\F_iw[11]~39_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[11]~q ),
	.prn(vcc));
defparam \D_iw[11] .is_wysiwyg = "true";
defparam \D_iw[11] .power_up = "low";

cyclone10lp_lcell_comb \F_iw[13]~40 (
	.dataa(src1_valid1),
	.datab(src1_valid2),
	.datac(q_a_13),
	.datad(av_readdata_pre_131),
	.cin(gnd),
	.combout(\F_iw[13]~40_combout ),
	.cout());
defparam \F_iw[13]~40 .lut_mask = 16'hFFFE;
defparam \F_iw[13]~40 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[13]~41 (
	.dataa(\F_iw[13]~40_combout ),
	.datab(src1_valid),
	.datac(av_readdata_pre_132),
	.datad(\D_iw[26]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[13]~41_combout ),
	.cout());
defparam \F_iw[13]~41 .lut_mask = 16'hFEFF;
defparam \F_iw[13]~41 .sum_lutc_input = "datac";

dffeas \D_iw[13] (
	.clk(clk_clk),
	.d(\F_iw[13]~41_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[13]~q ),
	.prn(vcc));
defparam \D_iw[13] .is_wysiwyg = "true";
defparam \D_iw[13] .power_up = "low";

cyclone10lp_lcell_comb \F_iw[16]~42 (
	.dataa(src1_valid1),
	.datab(src1_valid2),
	.datac(q_a_16),
	.datad(av_readdata_pre_161),
	.cin(gnd),
	.combout(\F_iw[16]~42_combout ),
	.cout());
defparam \F_iw[16]~42 .lut_mask = 16'hFFFE;
defparam \F_iw[16]~42 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[16]~43 (
	.dataa(\F_iw[16]~42_combout ),
	.datab(src1_valid),
	.datac(av_readdata_pre_16),
	.datad(\D_iw[26]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[16]~43_combout ),
	.cout());
defparam \F_iw[16]~43 .lut_mask = 16'hFEFF;
defparam \F_iw[16]~43 .sum_lutc_input = "datac";

dffeas \D_iw[16] (
	.clk(clk_clk),
	.d(\F_iw[16]~43_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[16]~q ),
	.prn(vcc));
defparam \D_iw[16] .is_wysiwyg = "true";
defparam \D_iw[16] .power_up = "low";

cyclone10lp_lcell_comb \F_iw[12]~44 (
	.dataa(src1_valid1),
	.datab(src1_valid2),
	.datac(q_a_12),
	.datad(av_readdata_pre_121),
	.cin(gnd),
	.combout(\F_iw[12]~44_combout ),
	.cout());
defparam \F_iw[12]~44 .lut_mask = 16'hFFFE;
defparam \F_iw[12]~44 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[12]~45 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[12]~44_combout ),
	.datac(src1_valid),
	.datad(av_readdata_pre_122),
	.cin(gnd),
	.combout(\F_iw[12]~45_combout ),
	.cout());
defparam \F_iw[12]~45 .lut_mask = 16'hFFFE;
defparam \F_iw[12]~45 .sum_lutc_input = "datac";

dffeas \D_iw[12] (
	.clk(clk_clk),
	.d(\F_iw[12]~45_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[12]~q ),
	.prn(vcc));
defparam \D_iw[12] .is_wysiwyg = "true";
defparam \D_iw[12] .power_up = "low";

cyclone10lp_lcell_comb \Equal62~7 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~7_combout ),
	.cout());
defparam \Equal62~7 .lut_mask = 16'hFF7F;
defparam \Equal62~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal62~9 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~9_combout ),
	.cout());
defparam \Equal62~9 .lut_mask = 16'hFFF7;
defparam \Equal62~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal62~10 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~10_combout ),
	.cout());
defparam \Equal62~10 .lut_mask = 16'hFFFB;
defparam \Equal62~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_shift_rot~0 (
	.dataa(\D_op_opx_rsv63~0_combout ),
	.datab(\Equal62~7_combout ),
	.datac(\Equal62~9_combout ),
	.datad(\Equal62~10_combout ),
	.cin(gnd),
	.combout(\D_ctrl_shift_rot~0_combout ),
	.cout());
defparam \D_ctrl_shift_rot~0 .lut_mask = 16'hFFFE;
defparam \D_ctrl_shift_rot~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_shift_logical~0 (
	.dataa(\D_iw[12]~q ),
	.datab(gnd),
	.datac(\D_iw[13]~q ),
	.datad(\D_iw[16]~q ),
	.cin(gnd),
	.combout(\D_ctrl_shift_logical~0_combout ),
	.cout());
defparam \D_ctrl_shift_logical~0 .lut_mask = 16'hAFFF;
defparam \D_ctrl_shift_logical~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_shift_rot~1 (
	.dataa(\D_ctrl_shift_logical~0_combout ),
	.datab(\Equal62~7_combout ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_shift_rot~1_combout ),
	.cout());
defparam \D_ctrl_shift_rot~1 .lut_mask = 16'hACFF;
defparam \D_ctrl_shift_rot~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal62~14 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~14_combout ),
	.cout());
defparam \Equal62~14 .lut_mask = 16'hFFBF;
defparam \Equal62~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_shift_rot~2 (
	.dataa(\D_ctrl_shift_rot~1_combout ),
	.datab(\Equal62~14_combout ),
	.datac(\D_iw[14]~q ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_ctrl_shift_rot~2_combout ),
	.cout());
defparam \D_ctrl_shift_rot~2 .lut_mask = 16'hFEFF;
defparam \D_ctrl_shift_rot~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_shift_rot~3 (
	.dataa(\Equal0~9_combout ),
	.datab(\D_ctrl_shift_rot~0_combout ),
	.datac(\D_ctrl_shift_rot~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_shift_rot~3_combout ),
	.cout());
defparam \D_ctrl_shift_rot~3 .lut_mask = 16'hFEFE;
defparam \D_ctrl_shift_rot~3 .sum_lutc_input = "datac";

dffeas R_ctrl_shift_rot(
	.clk(clk_clk),
	.d(\D_ctrl_shift_rot~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_shift_rot~q ),
	.prn(vcc));
defparam R_ctrl_shift_rot.is_wysiwyg = "true";
defparam R_ctrl_shift_rot.power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_cnt[0]~5 (
	.dataa(\E_shift_rot_cnt[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\E_shift_rot_cnt[0]~5_combout ),
	.cout(\E_shift_rot_cnt[0]~6 ));
defparam \E_shift_rot_cnt[0]~5 .lut_mask = 16'h55AA;
defparam \E_shift_rot_cnt[0]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_hi_imm16~0 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[4]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_hi_imm16~0_combout ),
	.cout());
defparam \D_ctrl_hi_imm16~0 .lut_mask = 16'hFFF7;
defparam \D_ctrl_hi_imm16~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_hi_imm16~1 (
	.dataa(\D_iw[2]~q ),
	.datab(\D_iw[5]~q ),
	.datac(\D_ctrl_hi_imm16~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_hi_imm16~1_combout ),
	.cout());
defparam \D_ctrl_hi_imm16~1 .lut_mask = 16'hFEFE;
defparam \D_ctrl_hi_imm16~1 .sum_lutc_input = "datac";

dffeas R_ctrl_hi_imm16(
	.clk(clk_clk),
	.d(\D_ctrl_hi_imm16~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_hi_imm16~q ),
	.prn(vcc));
defparam R_ctrl_hi_imm16.is_wysiwyg = "true";
defparam R_ctrl_hi_imm16.power_up = "low";

cyclone10lp_lcell_comb \D_ctrl_alu_force_xor~14 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[2]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[0]~q ),
	.cin(gnd),
	.combout(\D_ctrl_alu_force_xor~14_combout ),
	.cout());
defparam \D_ctrl_alu_force_xor~14 .lut_mask = 16'hF6FF;
defparam \D_ctrl_alu_force_xor~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal0~14 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~14_combout ),
	.cout());
defparam \Equal0~14 .lut_mask = 16'hFFFE;
defparam \Equal0~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal0~15 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~15_combout ),
	.cout());
defparam \Equal0~15 .lut_mask = 16'hFFFD;
defparam \Equal0~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_implicit_dst_eretaddr~3 (
	.dataa(\D_iw[5]~q ),
	.datab(\D_ctrl_alu_force_xor~14_combout ),
	.datac(\Equal0~14_combout ),
	.datad(\Equal0~15_combout ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~3_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~3 .lut_mask = 16'h7FFF;
defparam \D_ctrl_implicit_dst_eretaddr~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal62~5 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~5_combout ),
	.cout());
defparam \Equal62~5 .lut_mask = 16'hFEFF;
defparam \Equal62~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal62~12 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~12_combout ),
	.cout());
defparam \Equal62~12 .lut_mask = 16'hFDFF;
defparam \Equal62~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_force_src2_zero~0 (
	.dataa(\D_iw[15]~q ),
	.datab(\Equal62~5_combout ),
	.datac(\Equal62~12_combout ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~0_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_force_src2_zero~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal62~3 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~3_combout ),
	.cout());
defparam \Equal62~3 .lut_mask = 16'hEFFF;
defparam \Equal62~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_force_src2_zero~1 (
	.dataa(\Equal0~9_combout ),
	.datab(\D_ctrl_force_src2_zero~0_combout ),
	.datac(\Equal62~3_combout ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~1_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~1 .lut_mask = 16'hFEFF;
defparam \D_ctrl_force_src2_zero~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal62~4 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~4_combout ),
	.cout());
defparam \Equal62~4 .lut_mask = 16'hBFFF;
defparam \Equal62~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_uncond_cti_non_br~1 (
	.dataa(\D_iw[15]~q ),
	.datab(gnd),
	.datac(\Equal0~9_combout ),
	.datad(\Equal62~4_combout ),
	.cin(gnd),
	.combout(\D_ctrl_uncond_cti_non_br~1_combout ),
	.cout());
defparam \D_ctrl_uncond_cti_non_br~1 .lut_mask = 16'hAFFF;
defparam \D_ctrl_uncond_cti_non_br~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal0~12 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~12_combout ),
	.cout());
defparam \Equal0~12 .lut_mask = 16'hDFFF;
defparam \Equal0~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal62~6 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~6_combout ),
	.cout());
defparam \Equal62~6 .lut_mask = 16'hFFEF;
defparam \Equal62~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_exception~4 (
	.dataa(gnd),
	.datab(\Equal62~6_combout ),
	.datac(\Equal62~7_combout ),
	.datad(\D_op_cmpge~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~4_combout ),
	.cout());
defparam \D_ctrl_exception~4 .lut_mask = 16'h3FFF;
defparam \D_ctrl_exception~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal62~8 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~8_combout ),
	.cout());
defparam \Equal62~8 .lut_mask = 16'hDFFF;
defparam \Equal62~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal0~5 (
	.dataa(\D_iw[4]~q ),
	.datab(\D_iw[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal0~5_combout ),
	.cout());
defparam \Equal0~5 .lut_mask = 16'hEEEE;
defparam \Equal0~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_op_opx_rsv17~0 (
	.dataa(\Equal0~4_combout ),
	.datab(\Equal0~5_combout ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_op_opx_rsv17~0_combout ),
	.cout());
defparam \D_op_opx_rsv17~0 .lut_mask = 16'hFEFF;
defparam \D_op_opx_rsv17~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_exception~5 (
	.dataa(gnd),
	.datab(\Equal62~4_combout ),
	.datac(\Equal62~8_combout ),
	.datad(\D_op_opx_rsv17~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~5_combout ),
	.cout());
defparam \D_ctrl_exception~5 .lut_mask = 16'h3FFF;
defparam \D_ctrl_exception~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal62~0 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~0_combout ),
	.cout());
defparam \Equal62~0 .lut_mask = 16'h7FFF;
defparam \Equal62~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal62~2 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~2_combout ),
	.cout());
defparam \Equal62~2 .lut_mask = 16'hFBFF;
defparam \Equal62~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_op_opx_rsv00~0 (
	.dataa(\Equal0~4_combout ),
	.datab(\Equal0~5_combout ),
	.datac(\D_iw[14]~q ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_op_opx_rsv00~0_combout ),
	.cout());
defparam \D_op_opx_rsv00~0 .lut_mask = 16'hEFFF;
defparam \D_op_opx_rsv00~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_exception~6 (
	.dataa(gnd),
	.datab(\Equal62~0_combout ),
	.datac(\Equal62~2_combout ),
	.datad(\D_op_opx_rsv00~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~6_combout ),
	.cout());
defparam \D_ctrl_exception~6 .lut_mask = 16'h3FFF;
defparam \D_ctrl_exception~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_exception~7 (
	.dataa(gnd),
	.datab(\Equal62~9_combout ),
	.datac(\Equal62~10_combout ),
	.datad(\D_op_opx_rsv00~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~7_combout ),
	.cout());
defparam \D_ctrl_exception~7 .lut_mask = 16'h3FFF;
defparam \D_ctrl_exception~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_exception~8 (
	.dataa(\D_ctrl_exception~4_combout ),
	.datab(\D_ctrl_exception~5_combout ),
	.datac(\D_ctrl_exception~6_combout ),
	.datad(\D_ctrl_exception~7_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~8_combout ),
	.cout());
defparam \D_ctrl_exception~8 .lut_mask = 16'hFFFE;
defparam \D_ctrl_exception~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_exception~9 (
	.dataa(gnd),
	.datab(\Equal62~9_combout ),
	.datac(\Equal62~3_combout ),
	.datad(\D_op_opx_rsv17~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~9_combout ),
	.cout());
defparam \D_ctrl_exception~9 .lut_mask = 16'h3FFF;
defparam \D_ctrl_exception~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_exception~10 (
	.dataa(\D_ctrl_exception~9_combout ),
	.datab(\Equal62~9_combout ),
	.datac(\Equal62~10_combout ),
	.datad(\D_op_cmpge~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~10_combout ),
	.cout());
defparam \D_ctrl_exception~10 .lut_mask = 16'hBFFF;
defparam \D_ctrl_exception~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal62~1 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~1_combout ),
	.cout());
defparam \Equal62~1 .lut_mask = 16'hF7FF;
defparam \Equal62~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_exception~11 (
	.dataa(\Equal62~4_combout ),
	.datab(\Equal62~1_combout ),
	.datac(\Equal0~9_combout ),
	.datad(\D_op_opx_rsv63~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~11_combout ),
	.cout());
defparam \D_ctrl_exception~11 .lut_mask = 16'h7FFF;
defparam \D_ctrl_exception~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal62~11 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~11_combout ),
	.cout());
defparam \Equal62~11 .lut_mask = 16'hFFFE;
defparam \Equal62~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_exception~12 (
	.dataa(\D_iw[14]~q ),
	.datab(\D_iw[15]~q ),
	.datac(\Equal0~9_combout ),
	.datad(\Equal62~11_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~12_combout ),
	.cout());
defparam \D_ctrl_exception~12 .lut_mask = 16'h7FFF;
defparam \D_ctrl_exception~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal62~13 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~13_combout ),
	.cout());
defparam \Equal62~13 .lut_mask = 16'hFFFD;
defparam \Equal62~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_exception~13 (
	.dataa(\Equal62~12_combout ),
	.datab(\Equal62~13_combout ),
	.datac(\Equal0~9_combout ),
	.datad(\D_op_opx_rsv63~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~13_combout ),
	.cout());
defparam \D_ctrl_exception~13 .lut_mask = 16'h7FFF;
defparam \D_ctrl_exception~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal0~10 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~10_combout ),
	.cout());
defparam \Equal0~10 .lut_mask = 16'hFDFF;
defparam \Equal0~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_exception~14 (
	.dataa(\D_ctrl_exception~13_combout ),
	.datab(\D_op_opx_rsv17~0_combout ),
	.datac(\Equal62~10_combout ),
	.datad(\Equal0~10_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~14_combout ),
	.cout());
defparam \D_ctrl_exception~14 .lut_mask = 16'hBFFF;
defparam \D_ctrl_exception~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_exception~15 (
	.dataa(\D_ctrl_exception~10_combout ),
	.datab(\D_ctrl_exception~11_combout ),
	.datac(\D_ctrl_exception~12_combout ),
	.datad(\D_ctrl_exception~14_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~15_combout ),
	.cout());
defparam \D_ctrl_exception~15 .lut_mask = 16'hFFFE;
defparam \D_ctrl_exception~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal0~11 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~11_combout ),
	.cout());
defparam \Equal0~11 .lut_mask = 16'hBFFF;
defparam \Equal0~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal0~7 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~7_combout ),
	.cout());
defparam \Equal0~7 .lut_mask = 16'h7FFF;
defparam \Equal0~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_jmp_direct~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\D_iw[4]~q ),
	.datad(\D_iw[5]~q ),
	.cin(gnd),
	.combout(\D_ctrl_jmp_direct~0_combout ),
	.cout());
defparam \D_ctrl_jmp_direct~0 .lut_mask = 16'h0FFF;
defparam \D_ctrl_jmp_direct~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_retaddr~0 (
	.dataa(\D_iw[15]~q ),
	.datab(\Equal62~8_combout ),
	.datac(\Equal62~3_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~0_combout ),
	.cout());
defparam \D_ctrl_retaddr~0 .lut_mask = 16'hFEFE;
defparam \D_ctrl_retaddr~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_retaddr~1 (
	.dataa(\Equal62~5_combout ),
	.datab(\Equal62~12_combout ),
	.datac(gnd),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~1_combout ),
	.cout());
defparam \D_ctrl_retaddr~1 .lut_mask = 16'hEEFF;
defparam \D_ctrl_retaddr~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_retaddr~2 (
	.dataa(\Equal0~9_combout ),
	.datab(\D_iw[14]~q ),
	.datac(\D_ctrl_retaddr~0_combout ),
	.datad(\D_ctrl_retaddr~1_combout ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~2_combout ),
	.cout());
defparam \D_ctrl_retaddr~2 .lut_mask = 16'hFFFE;
defparam \D_ctrl_retaddr~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_force_src2_zero~2 (
	.dataa(\Equal0~11_combout ),
	.datab(\Equal0~7_combout ),
	.datac(\D_ctrl_jmp_direct~0_combout ),
	.datad(\D_ctrl_retaddr~2_combout ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~2_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~2 .lut_mask = 16'h7FFF;
defparam \D_ctrl_force_src2_zero~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal0~21 (
	.dataa(\Equal0~4_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\D_iw[5]~q ),
	.cin(gnd),
	.combout(\Equal0~21_combout ),
	.cout());
defparam \Equal0~21 .lut_mask = 16'hAAFF;
defparam \Equal0~21 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_force_src2_zero~3 (
	.dataa(\D_ctrl_exception~8_combout ),
	.datab(\D_ctrl_exception~15_combout ),
	.datac(\D_ctrl_force_src2_zero~2_combout ),
	.datad(\Equal0~21_combout ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~3_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~3 .lut_mask = 16'hFEFF;
defparam \D_ctrl_force_src2_zero~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_force_src2_zero~4 (
	.dataa(\D_ctrl_force_src2_zero~1_combout ),
	.datab(\D_ctrl_uncond_cti_non_br~1_combout ),
	.datac(\Equal0~12_combout ),
	.datad(\D_ctrl_force_src2_zero~3_combout ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~4_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~4 .lut_mask = 16'hFFDF;
defparam \D_ctrl_force_src2_zero~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_force_src2_zero~5 (
	.dataa(\D_iw[4]~q ),
	.datab(\Equal0~11_combout ),
	.datac(\D_iw[5]~q ),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~5_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~5 .lut_mask = 16'hFFDE;
defparam \D_ctrl_force_src2_zero~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_force_src2_zero~6 (
	.dataa(\D_ctrl_implicit_dst_eretaddr~3_combout ),
	.datab(\D_ctrl_force_src2_zero~4_combout ),
	.datac(\D_iw[4]~q ),
	.datad(\D_ctrl_force_src2_zero~5_combout ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~6_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~6 .lut_mask = 16'hFFF7;
defparam \D_ctrl_force_src2_zero~6 .sum_lutc_input = "datac";

dffeas R_ctrl_force_src2_zero(
	.clk(clk_clk),
	.d(\D_ctrl_force_src2_zero~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_force_src2_zero~q ),
	.prn(vcc));
defparam R_ctrl_force_src2_zero.is_wysiwyg = "true";
defparam R_ctrl_force_src2_zero.power_up = "low";

cyclone10lp_lcell_comb \R_src2_lo[4]~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\R_ctrl_hi_imm16~q ),
	.datad(\R_ctrl_force_src2_zero~q ),
	.cin(gnd),
	.combout(\R_src2_lo[4]~3_combout ),
	.cout());
defparam \R_src2_lo[4]~3 .lut_mask = 16'h0FFF;
defparam \R_src2_lo[4]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[6]~58 (
	.dataa(src1_valid),
	.datab(src1_valid1),
	.datac(av_readdata_pre_6),
	.datad(av_readdata_pre_61),
	.cin(gnd),
	.combout(\F_iw[6]~58_combout ),
	.cout());
defparam \F_iw[6]~58 .lut_mask = 16'hFFFE;
defparam \F_iw[6]~58 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[6]~59 (
	.dataa(read_latency_shift_reg_01),
	.datab(mem_74_01),
	.datac(mem_56_01),
	.datad(q_a_6),
	.cin(gnd),
	.combout(\F_iw[6]~59_combout ),
	.cout());
defparam \F_iw[6]~59 .lut_mask = 16'hFFFE;
defparam \F_iw[6]~59 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[6]~60 (
	.dataa(\F_iw[6]~58_combout ),
	.datab(\F_iw[6]~59_combout ),
	.datac(src1_valid3),
	.datad(av_readdata_pre_62),
	.cin(gnd),
	.combout(\F_iw[6]~60_combout ),
	.cout());
defparam \F_iw[6]~60 .lut_mask = 16'hFFFE;
defparam \F_iw[6]~60 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[6]~61 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[6]~60_combout ),
	.datac(src1_valid4),
	.datad(av_readdata_pre_63),
	.cin(gnd),
	.combout(\F_iw[6]~61_combout ),
	.cout());
defparam \F_iw[6]~61 .lut_mask = 16'hFFFE;
defparam \F_iw[6]~61 .sum_lutc_input = "datac";

dffeas \D_iw[6] (
	.clk(clk_clk),
	.d(\F_iw[6]~61_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[6]~q ),
	.prn(vcc));
defparam \D_iw[6] .is_wysiwyg = "true";
defparam \D_iw[6] .power_up = "low";

cyclone10lp_lcell_comb \D_ctrl_implicit_dst_eretaddr~0 (
	.dataa(\D_iw[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~0_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~0 .lut_mask = 16'hAAFF;
defparam \D_ctrl_implicit_dst_eretaddr~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_unsigned_lo_imm16~2 (
	.dataa(\D_op_opx_rsv63~0_combout ),
	.datab(\Equal62~9_combout ),
	.datac(\Equal62~7_combout ),
	.datad(\D_ctrl_implicit_dst_eretaddr~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_unsigned_lo_imm16~2_combout ),
	.cout());
defparam \D_ctrl_unsigned_lo_imm16~2 .lut_mask = 16'hFEFF;
defparam \D_ctrl_unsigned_lo_imm16~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_unsigned_lo_imm16~5 (
	.dataa(\D_iw[4]~q ),
	.datab(\Equal0~4_combout ),
	.datac(\D_iw[5]~q ),
	.datad(\D_ctrl_unsigned_lo_imm16~2_combout ),
	.cin(gnd),
	.combout(\D_ctrl_unsigned_lo_imm16~5_combout ),
	.cout());
defparam \D_ctrl_unsigned_lo_imm16~5 .lut_mask = 16'hFFFE;
defparam \D_ctrl_unsigned_lo_imm16~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_b_is_dst~0 (
	.dataa(\D_iw[2]~q ),
	.datab(\D_iw[3]~q ),
	.datac(\D_iw[5]~q ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_b_is_dst~0_combout ),
	.cout());
defparam \D_ctrl_b_is_dst~0 .lut_mask = 16'h6996;
defparam \D_ctrl_b_is_dst~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_b_is_dst~1 (
	.dataa(\D_iw[2]~q ),
	.datab(\D_iw[3]~q ),
	.datac(\D_iw[5]~q ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_b_is_dst~1_combout ),
	.cout());
defparam \D_ctrl_b_is_dst~1 .lut_mask = 16'hFBFE;
defparam \D_ctrl_b_is_dst~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_b_is_dst~2 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[1]~q ),
	.datac(\D_ctrl_b_is_dst~0_combout ),
	.datad(\D_ctrl_b_is_dst~1_combout ),
	.cin(gnd),
	.combout(\D_ctrl_b_is_dst~2_combout ),
	.cout());
defparam \D_ctrl_b_is_dst~2 .lut_mask = 16'h96FF;
defparam \D_ctrl_b_is_dst~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal0~18 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~18_combout ),
	.cout());
defparam \Equal0~18 .lut_mask = 16'hFFDF;
defparam \Equal0~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_src2_use_imm~0 (
	.dataa(\D_ctrl_b_is_dst~2_combout ),
	.datab(\Equal0~18_combout ),
	.datac(\Equal0~15_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\R_src2_use_imm~0_combout ),
	.cout());
defparam \R_src2_use_imm~0 .lut_mask = 16'hFEFF;
defparam \R_src2_use_imm~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_ctrl_br_nxt~0 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[4]~q ),
	.datac(\D_iw[5]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\R_ctrl_br_nxt~0_combout ),
	.cout());
defparam \R_ctrl_br_nxt~0 .lut_mask = 16'hFFFE;
defparam \R_ctrl_br_nxt~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_ctrl_br_nxt~1 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[2]~q ),
	.datac(gnd),
	.datad(\R_ctrl_br_nxt~0_combout ),
	.cin(gnd),
	.combout(\R_ctrl_br_nxt~1_combout ),
	.cout());
defparam \R_ctrl_br_nxt~1 .lut_mask = 16'hEEFF;
defparam \R_ctrl_br_nxt~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_src2_use_imm~1 (
	.dataa(\D_ctrl_unsigned_lo_imm16~5_combout ),
	.datab(\R_src2_use_imm~0_combout ),
	.datac(\R_ctrl_br_nxt~1_combout ),
	.datad(\R_valid~q ),
	.cin(gnd),
	.combout(\R_src2_use_imm~1_combout ),
	.cout());
defparam \R_src2_use_imm~1 .lut_mask = 16'hFFFE;
defparam \R_src2_use_imm~1 .sum_lutc_input = "datac";

dffeas R_src2_use_imm(
	.clk(clk_clk),
	.d(\R_src2_use_imm~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_src2_use_imm~q ),
	.prn(vcc));
defparam R_src2_use_imm.is_wysiwyg = "true";
defparam R_src2_use_imm.power_up = "low";

cyclone10lp_lcell_comb \D_ctrl_src_imm5_shift_rot~0 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[15]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_src_imm5_shift_rot~0_combout ),
	.cout());
defparam \D_ctrl_src_imm5_shift_rot~0 .lut_mask = 16'hBBF3;
defparam \D_ctrl_src_imm5_shift_rot~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_src_imm5_shift_rot~1 (
	.dataa(\Equal0~9_combout ),
	.datab(\D_iw[12]~q ),
	.datac(\D_iw[13]~q ),
	.datad(\D_ctrl_src_imm5_shift_rot~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_src_imm5_shift_rot~1_combout ),
	.cout());
defparam \D_ctrl_src_imm5_shift_rot~1 .lut_mask = 16'hEFFF;
defparam \D_ctrl_src_imm5_shift_rot~1 .sum_lutc_input = "datac";

dffeas R_ctrl_src_imm5_shift_rot(
	.clk(clk_clk),
	.d(\D_ctrl_src_imm5_shift_rot~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_src_imm5_shift_rot~q ),
	.prn(vcc));
defparam R_ctrl_src_imm5_shift_rot.is_wysiwyg = "true";
defparam R_ctrl_src_imm5_shift_rot.power_up = "low";

cyclone10lp_lcell_comb \R_src2_lo~4 (
	.dataa(\R_src2_use_imm~q ),
	.datab(\R_ctrl_src_imm5_shift_rot~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\R_src2_lo~4_combout ),
	.cout());
defparam \R_src2_lo~4 .lut_mask = 16'hEEEE;
defparam \R_src2_lo~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_src2_lo[0]~9 (
	.dataa(\R_src2_lo[4]~3_combout ),
	.datab(\D_iw[6]~q ),
	.datac(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.datad(\R_src2_lo~4_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[0]~9_combout ),
	.cout());
defparam \R_src2_lo[0]~9 .lut_mask = 16'hFAFC;
defparam \R_src2_lo[0]~9 .sum_lutc_input = "datac";

dffeas \E_src2[0] (
	.clk(clk_clk),
	.d(\R_src2_lo[0]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[0]~q ),
	.prn(vcc));
defparam \E_src2[0] .is_wysiwyg = "true";
defparam \E_src2[0] .power_up = "low";

dffeas \E_shift_rot_cnt[0] (
	.clk(clk_clk),
	.d(\E_shift_rot_cnt[0]~5_combout ),
	.asdata(\E_src2[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[0]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[0] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[0] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_cnt[1]~7 (
	.dataa(\E_shift_rot_cnt[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\E_shift_rot_cnt[0]~6 ),
	.combout(\E_shift_rot_cnt[1]~7_combout ),
	.cout(\E_shift_rot_cnt[1]~8 ));
defparam \E_shift_rot_cnt[1]~7 .lut_mask = 16'h5A5F;
defparam \E_shift_rot_cnt[1]~7 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \F_iw[7]~54 (
	.dataa(src1_valid),
	.datab(src1_valid1),
	.datac(av_readdata_pre_7),
	.datad(av_readdata_pre_71),
	.cin(gnd),
	.combout(\F_iw[7]~54_combout ),
	.cout());
defparam \F_iw[7]~54 .lut_mask = 16'hFFFE;
defparam \F_iw[7]~54 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[7]~55 (
	.dataa(read_latency_shift_reg_01),
	.datab(mem_74_01),
	.datac(mem_56_01),
	.datad(q_a_7),
	.cin(gnd),
	.combout(\F_iw[7]~55_combout ),
	.cout());
defparam \F_iw[7]~55 .lut_mask = 16'hFFFE;
defparam \F_iw[7]~55 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[7]~56 (
	.dataa(\F_iw[7]~54_combout ),
	.datab(\F_iw[7]~55_combout ),
	.datac(src1_valid3),
	.datad(av_readdata_pre_72),
	.cin(gnd),
	.combout(\F_iw[7]~56_combout ),
	.cout());
defparam \F_iw[7]~56 .lut_mask = 16'hFFFE;
defparam \F_iw[7]~56 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[7]~57 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[7]~56_combout ),
	.datac(src1_valid4),
	.datad(av_readdata_pre_73),
	.cin(gnd),
	.combout(\F_iw[7]~57_combout ),
	.cout());
defparam \F_iw[7]~57 .lut_mask = 16'hFFFE;
defparam \F_iw[7]~57 .sum_lutc_input = "datac";

dffeas \D_iw[7] (
	.clk(clk_clk),
	.d(\F_iw[7]~57_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[7]~q ),
	.prn(vcc));
defparam \D_iw[7] .is_wysiwyg = "true";
defparam \D_iw[7] .power_up = "low";

cyclone10lp_lcell_comb \R_src2_lo[1]~8 (
	.dataa(\R_src2_lo[4]~3_combout ),
	.datab(\D_iw[7]~q ),
	.datac(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.datad(\R_src2_lo~4_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[1]~8_combout ),
	.cout());
defparam \R_src2_lo[1]~8 .lut_mask = 16'hFAFC;
defparam \R_src2_lo[1]~8 .sum_lutc_input = "datac";

dffeas \E_src2[1] (
	.clk(clk_clk),
	.d(\R_src2_lo[1]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[1]~q ),
	.prn(vcc));
defparam \E_src2[1] .is_wysiwyg = "true";
defparam \E_src2[1] .power_up = "low";

dffeas \E_shift_rot_cnt[1] (
	.clk(clk_clk),
	.d(\E_shift_rot_cnt[1]~7_combout ),
	.asdata(\E_src2[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[1]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[1] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[1] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_cnt[2]~9 (
	.dataa(\E_shift_rot_cnt[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\E_shift_rot_cnt[1]~8 ),
	.combout(\E_shift_rot_cnt[2]~9_combout ),
	.cout(\E_shift_rot_cnt[2]~10 ));
defparam \E_shift_rot_cnt[2]~9 .lut_mask = 16'h5AAF;
defparam \E_shift_rot_cnt[2]~9 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \F_iw[8]~51 (
	.dataa(src1_valid),
	.datab(src1_valid1),
	.datac(av_readdata_pre_8),
	.datad(av_readdata_pre_81),
	.cin(gnd),
	.combout(\F_iw[8]~51_combout ),
	.cout());
defparam \F_iw[8]~51 .lut_mask = 16'hFFFE;
defparam \F_iw[8]~51 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[8]~52 (
	.dataa(src1_valid2),
	.datab(src1_valid4),
	.datac(av_readdata_pre_82),
	.datad(q_a_8),
	.cin(gnd),
	.combout(\F_iw[8]~52_combout ),
	.cout());
defparam \F_iw[8]~52 .lut_mask = 16'hFFFE;
defparam \F_iw[8]~52 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[8]~53 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[8]~51_combout ),
	.datac(\F_iw[8]~52_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\F_iw[8]~53_combout ),
	.cout());
defparam \F_iw[8]~53 .lut_mask = 16'hFEFE;
defparam \F_iw[8]~53 .sum_lutc_input = "datac";

dffeas \D_iw[8] (
	.clk(clk_clk),
	.d(\F_iw[8]~53_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[8]~q ),
	.prn(vcc));
defparam \D_iw[8] .is_wysiwyg = "true";
defparam \D_iw[8] .power_up = "low";

cyclone10lp_lcell_comb \R_src2_lo[2]~7 (
	.dataa(\R_src2_lo[4]~3_combout ),
	.datab(\D_iw[8]~q ),
	.datac(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.datad(\R_src2_lo~4_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[2]~7_combout ),
	.cout());
defparam \R_src2_lo[2]~7 .lut_mask = 16'hFAFC;
defparam \R_src2_lo[2]~7 .sum_lutc_input = "datac";

dffeas \E_src2[2] (
	.clk(clk_clk),
	.d(\R_src2_lo[2]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[2]~q ),
	.prn(vcc));
defparam \E_src2[2] .is_wysiwyg = "true";
defparam \E_src2[2] .power_up = "low";

dffeas \E_shift_rot_cnt[2] (
	.clk(clk_clk),
	.d(\E_shift_rot_cnt[2]~9_combout ),
	.asdata(\E_src2[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[2]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[2] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[2] .power_up = "low";

cyclone10lp_lcell_comb \E_stall~0 (
	.dataa(\E_new_inst~q ),
	.datab(\E_shift_rot_cnt[0]~q ),
	.datac(\E_shift_rot_cnt[1]~q ),
	.datad(\E_shift_rot_cnt[2]~q ),
	.cin(gnd),
	.combout(\E_stall~0_combout ),
	.cout());
defparam \E_stall~0 .lut_mask = 16'hFFFE;
defparam \E_stall~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_shift_rot_cnt[3]~11 (
	.dataa(\E_shift_rot_cnt[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\E_shift_rot_cnt[2]~10 ),
	.combout(\E_shift_rot_cnt[3]~11_combout ),
	.cout(\E_shift_rot_cnt[3]~12 ));
defparam \E_shift_rot_cnt[3]~11 .lut_mask = 16'h5A5F;
defparam \E_shift_rot_cnt[3]~11 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \F_iw[9]~48 (
	.dataa(src1_valid),
	.datab(src1_valid1),
	.datac(av_readdata_pre_9),
	.datad(av_readdata_pre_91),
	.cin(gnd),
	.combout(\F_iw[9]~48_combout ),
	.cout());
defparam \F_iw[9]~48 .lut_mask = 16'hFFFE;
defparam \F_iw[9]~48 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[9]~49 (
	.dataa(src1_valid2),
	.datab(src1_valid4),
	.datac(av_readdata_pre_92),
	.datad(q_a_9),
	.cin(gnd),
	.combout(\F_iw[9]~49_combout ),
	.cout());
defparam \F_iw[9]~49 .lut_mask = 16'hFFFE;
defparam \F_iw[9]~49 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[9]~50 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[9]~48_combout ),
	.datac(\F_iw[9]~49_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\F_iw[9]~50_combout ),
	.cout());
defparam \F_iw[9]~50 .lut_mask = 16'hFEFE;
defparam \F_iw[9]~50 .sum_lutc_input = "datac";

dffeas \D_iw[9] (
	.clk(clk_clk),
	.d(\F_iw[9]~50_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[9]~q ),
	.prn(vcc));
defparam \D_iw[9] .is_wysiwyg = "true";
defparam \D_iw[9] .power_up = "low";

cyclone10lp_lcell_comb \R_src2_lo[3]~6 (
	.dataa(\R_src2_lo[4]~3_combout ),
	.datab(\D_iw[9]~q ),
	.datac(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.datad(\R_src2_lo~4_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[3]~6_combout ),
	.cout());
defparam \R_src2_lo[3]~6 .lut_mask = 16'hFAFC;
defparam \R_src2_lo[3]~6 .sum_lutc_input = "datac";

dffeas \E_src2[3] (
	.clk(clk_clk),
	.d(\R_src2_lo[3]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[3]~q ),
	.prn(vcc));
defparam \E_src2[3] .is_wysiwyg = "true";
defparam \E_src2[3] .power_up = "low";

dffeas \E_shift_rot_cnt[3] (
	.clk(clk_clk),
	.d(\E_shift_rot_cnt[3]~11_combout ),
	.asdata(\E_src2[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[3]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[3] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[3] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_cnt[4]~13 (
	.dataa(\E_shift_rot_cnt[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\E_shift_rot_cnt[3]~12 ),
	.combout(\E_shift_rot_cnt[4]~13_combout ),
	.cout());
defparam \E_shift_rot_cnt[4]~13 .lut_mask = 16'h5A5A;
defparam \E_shift_rot_cnt[4]~13 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \F_iw[10]~46 (
	.dataa(src1_valid1),
	.datab(src1_valid2),
	.datac(q_a_10),
	.datad(av_readdata_pre_10),
	.cin(gnd),
	.combout(\F_iw[10]~46_combout ),
	.cout());
defparam \F_iw[10]~46 .lut_mask = 16'hFFFE;
defparam \F_iw[10]~46 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[10]~47 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[10]~46_combout ),
	.datac(src1_valid),
	.datad(av_readdata_pre_101),
	.cin(gnd),
	.combout(\F_iw[10]~47_combout ),
	.cout());
defparam \F_iw[10]~47 .lut_mask = 16'hFFFE;
defparam \F_iw[10]~47 .sum_lutc_input = "datac";

dffeas \D_iw[10] (
	.clk(clk_clk),
	.d(\F_iw[10]~47_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[10]~q ),
	.prn(vcc));
defparam \D_iw[10] .is_wysiwyg = "true";
defparam \D_iw[10] .power_up = "low";

cyclone10lp_lcell_comb \R_src2_lo[4]~5 (
	.dataa(\R_src2_lo[4]~3_combout ),
	.datab(\D_iw[10]~q ),
	.datac(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.datad(\R_src2_lo~4_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[4]~5_combout ),
	.cout());
defparam \R_src2_lo[4]~5 .lut_mask = 16'hFAFC;
defparam \R_src2_lo[4]~5 .sum_lutc_input = "datac";

dffeas \E_src2[4] (
	.clk(clk_clk),
	.d(\R_src2_lo[4]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[4]~q ),
	.prn(vcc));
defparam \E_src2[4] .is_wysiwyg = "true";
defparam \E_src2[4] .power_up = "low";

dffeas \E_shift_rot_cnt[4] (
	.clk(clk_clk),
	.d(\E_shift_rot_cnt[4]~13_combout ),
	.asdata(\E_src2[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[4]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[4] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[4] .power_up = "low";

cyclone10lp_lcell_comb \E_stall~1 (
	.dataa(\E_shift_rot_cnt[3]~q ),
	.datab(\E_shift_rot_cnt[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\E_stall~1_combout ),
	.cout());
defparam \E_stall~1 .lut_mask = 16'hEEEE;
defparam \E_stall~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_stall~2 (
	.dataa(\R_ctrl_shift_rot~q ),
	.datab(\E_valid_from_R~q ),
	.datac(\E_stall~0_combout ),
	.datad(\E_stall~1_combout ),
	.cin(gnd),
	.combout(\E_stall~2_combout ),
	.cout());
defparam \E_stall~2 .lut_mask = 16'hFFFE;
defparam \E_stall~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_ld_signed~0 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[4]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_ld_signed~0_combout ),
	.cout());
defparam \D_ctrl_ld_signed~0 .lut_mask = 16'hEFFF;
defparam \D_ctrl_ld_signed~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_ld~2 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[2]~q ),
	.datac(\D_iw[4]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_ld~2_combout ),
	.cout());
defparam \D_ctrl_ld~2 .lut_mask = 16'hBFBF;
defparam \D_ctrl_ld~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_ld~3 (
	.dataa(\D_iw[2]~q ),
	.datab(\D_ctrl_ld_signed~0_combout ),
	.datac(\D_iw[0]~q ),
	.datad(\D_ctrl_ld~2_combout ),
	.cin(gnd),
	.combout(\D_ctrl_ld~3_combout ),
	.cout());
defparam \D_ctrl_ld~3 .lut_mask = 16'hFFFE;
defparam \D_ctrl_ld~3 .sum_lutc_input = "datac";

dffeas R_ctrl_ld(
	.clk(clk_clk),
	.d(\D_ctrl_ld~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_ld~q ),
	.prn(vcc));
defparam R_ctrl_ld.is_wysiwyg = "true";
defparam R_ctrl_ld.power_up = "low";

dffeas av_ld_waiting_for_data(
	.clk(clk_clk),
	.d(\av_ld_waiting_for_data_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_waiting_for_data~q ),
	.prn(vcc));
defparam av_ld_waiting_for_data.is_wysiwyg = "true";
defparam av_ld_waiting_for_data.power_up = "low";

cyclone10lp_lcell_comb \av_ld_aligning_data_nxt~0 (
	.dataa(d_read1),
	.datab(gnd),
	.datac(WideOr1),
	.datad(WideOr11),
	.cin(gnd),
	.combout(\av_ld_aligning_data_nxt~0_combout ),
	.cout());
defparam \av_ld_aligning_data_nxt~0 .lut_mask = 16'hAFFF;
defparam \av_ld_aligning_data_nxt~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_waiting_for_data_nxt~0 (
	.dataa(\E_new_inst~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\av_ld_waiting_for_data~q ),
	.datad(\av_ld_aligning_data_nxt~0_combout ),
	.cin(gnd),
	.combout(\av_ld_waiting_for_data_nxt~0_combout ),
	.cout());
defparam \av_ld_waiting_for_data_nxt~0 .lut_mask = 16'hACFF;
defparam \av_ld_waiting_for_data_nxt~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_mem16~0 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[2]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_mem16~0_combout ),
	.cout());
defparam \D_ctrl_mem16~0 .lut_mask = 16'hFFFE;
defparam \D_ctrl_mem16~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_align_cycle_nxt[0]~0 (
	.dataa(\av_ld_align_cycle[0]~q ),
	.datab(d_read1),
	.datac(WideOr1),
	.datad(WideOr11),
	.cin(gnd),
	.combout(\av_ld_align_cycle_nxt[0]~0_combout ),
	.cout());
defparam \av_ld_align_cycle_nxt[0]~0 .lut_mask = 16'hFFF7;
defparam \av_ld_align_cycle_nxt[0]~0 .sum_lutc_input = "datac";

dffeas \av_ld_align_cycle[0] (
	.clk(clk_clk),
	.d(\av_ld_align_cycle_nxt[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_align_cycle[0]~q ),
	.prn(vcc));
defparam \av_ld_align_cycle[0] .is_wysiwyg = "true";
defparam \av_ld_align_cycle[0] .power_up = "low";

cyclone10lp_lcell_comb \av_ld_align_cycle_nxt[1]~1 (
	.dataa(gnd),
	.datab(\av_ld_align_cycle[1]~q ),
	.datac(\av_ld_align_cycle[0]~q ),
	.datad(\av_ld_aligning_data_nxt~0_combout ),
	.cin(gnd),
	.combout(\av_ld_align_cycle_nxt[1]~1_combout ),
	.cout());
defparam \av_ld_align_cycle_nxt[1]~1 .lut_mask = 16'h3CFF;
defparam \av_ld_align_cycle_nxt[1]~1 .sum_lutc_input = "datac";

dffeas \av_ld_align_cycle[1] (
	.clk(clk_clk),
	.d(\av_ld_align_cycle_nxt[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_align_cycle[1]~q ),
	.prn(vcc));
defparam \av_ld_align_cycle[1] .is_wysiwyg = "true";
defparam \av_ld_align_cycle[1] .power_up = "low";

cyclone10lp_lcell_comb \av_ld_aligning_data_nxt~1 (
	.dataa(\D_ctrl_mem16~0_combout ),
	.datab(\D_iw[4]~q ),
	.datac(\av_ld_align_cycle[0]~q ),
	.datad(\av_ld_align_cycle[1]~q ),
	.cin(gnd),
	.combout(\av_ld_aligning_data_nxt~1_combout ),
	.cout());
defparam \av_ld_aligning_data_nxt~1 .lut_mask = 16'h96FF;
defparam \av_ld_aligning_data_nxt~1 .sum_lutc_input = "datac";

dffeas av_ld_aligning_data(
	.clk(clk_clk),
	.d(\av_ld_aligning_data_nxt~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_aligning_data~q ),
	.prn(vcc));
defparam av_ld_aligning_data.is_wysiwyg = "true";
defparam av_ld_aligning_data.power_up = "low";

cyclone10lp_lcell_comb \D_ctrl_mem32~0 (
	.dataa(\D_iw[4]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[2]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_mem32~0_combout ),
	.cout());
defparam \D_ctrl_mem32~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_mem32~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \av_ld_aligning_data_nxt~2 (
	.dataa(\av_ld_aligning_data_nxt~1_combout ),
	.datab(\av_ld_aligning_data~q ),
	.datac(\av_ld_aligning_data_nxt~0_combout ),
	.datad(\D_ctrl_mem32~0_combout ),
	.cin(gnd),
	.combout(\av_ld_aligning_data_nxt~2_combout ),
	.cout());
defparam \av_ld_aligning_data_nxt~2 .lut_mask = 16'hB8FF;
defparam \av_ld_aligning_data_nxt~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_stall~3 (
	.dataa(\E_valid_from_R~q ),
	.datab(\av_ld_waiting_for_data_nxt~0_combout ),
	.datac(\av_ld_aligning_data_nxt~2_combout ),
	.datad(\D_ctrl_mem32~0_combout ),
	.cin(gnd),
	.combout(\E_stall~3_combout ),
	.cout());
defparam \E_stall~3 .lut_mask = 16'hFEFF;
defparam \E_stall~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_stall~4 (
	.dataa(\E_stall~2_combout ),
	.datab(\R_ctrl_ld~q ),
	.datac(\E_new_inst~q ),
	.datad(\E_stall~3_combout ),
	.cin(gnd),
	.combout(\E_stall~4_combout ),
	.cout());
defparam \E_stall~4 .lut_mask = 16'hFFFE;
defparam \E_stall~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_valid_from_R~0 (
	.dataa(\E_st_stall~combout ),
	.datab(\E_stall~4_combout ),
	.datac(\R_valid~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\E_valid_from_R~0_combout ),
	.cout());
defparam \E_valid_from_R~0 .lut_mask = 16'hFEFE;
defparam \E_valid_from_R~0 .sum_lutc_input = "datac";

dffeas E_valid_from_R(
	.clk(clk_clk),
	.d(\E_valid_from_R~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_valid_from_R~q ),
	.prn(vcc));
defparam E_valid_from_R.is_wysiwyg = "true";
defparam E_valid_from_R.power_up = "low";

cyclone10lp_lcell_comb \D_ctrl_jmp_direct~1 (
	.dataa(\D_ctrl_jmp_direct~0_combout ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[2]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_jmp_direct~1_combout ),
	.cout());
defparam \D_ctrl_jmp_direct~1 .lut_mask = 16'hBFFF;
defparam \D_ctrl_jmp_direct~1 .sum_lutc_input = "datac";

dffeas R_ctrl_jmp_direct(
	.clk(clk_clk),
	.d(\D_ctrl_jmp_direct~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_jmp_direct~q ),
	.prn(vcc));
defparam R_ctrl_jmp_direct.is_wysiwyg = "true";
defparam R_ctrl_jmp_direct.power_up = "low";

dffeas R_ctrl_br(
	.clk(clk_clk),
	.d(\R_ctrl_br_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_br~q ),
	.prn(vcc));
defparam R_ctrl_br.is_wysiwyg = "true";
defparam R_ctrl_br.power_up = "low";

cyclone10lp_lcell_comb \D_ctrl_retaddr~3 (
	.dataa(\Equal62~12_combout ),
	.datab(\Equal62~11_combout ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~3_combout ),
	.cout());
defparam \D_ctrl_retaddr~3 .lut_mask = 16'hEFFF;
defparam \D_ctrl_retaddr~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_retaddr~4 (
	.dataa(\D_ctrl_retaddr~3_combout ),
	.datab(\Equal62~5_combout ),
	.datac(\Equal62~6_combout ),
	.datad(\D_ctrl_implicit_dst_eretaddr~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~4_combout ),
	.cout());
defparam \D_ctrl_retaddr~4 .lut_mask = 16'hFEFF;
defparam \D_ctrl_retaddr~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_retaddr~5 (
	.dataa(\Equal0~9_combout ),
	.datab(\D_ctrl_retaddr~4_combout ),
	.datac(\D_ctrl_force_src2_zero~3_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~5_combout ),
	.cout());
defparam \D_ctrl_retaddr~5 .lut_mask = 16'hF7F7;
defparam \D_ctrl_retaddr~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal0~13 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~13_combout ),
	.cout());
defparam \Equal0~13 .lut_mask = 16'hFF7F;
defparam \Equal0~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_retaddr~6 (
	.dataa(\Equal0~12_combout ),
	.datab(\D_ctrl_implicit_dst_eretaddr~3_combout ),
	.datac(\Equal0~13_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~6_combout ),
	.cout());
defparam \D_ctrl_retaddr~6 .lut_mask = 16'hFDFE;
defparam \D_ctrl_retaddr~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_retaddr~7 (
	.dataa(\D_iw[5]~q ),
	.datab(\Equal0~11_combout ),
	.datac(\D_iw[4]~q ),
	.datad(\D_ctrl_retaddr~6_combout ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~7_combout ),
	.cout());
defparam \D_ctrl_retaddr~7 .lut_mask = 16'hFFBE;
defparam \D_ctrl_retaddr~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_retaddr~8 (
	.dataa(\Equal0~4_combout ),
	.datab(\D_ctrl_retaddr~5_combout ),
	.datac(\D_iw[4]~q ),
	.datad(\D_ctrl_retaddr~7_combout ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~8_combout ),
	.cout());
defparam \D_ctrl_retaddr~8 .lut_mask = 16'hBFFB;
defparam \D_ctrl_retaddr~8 .sum_lutc_input = "datac";

dffeas R_ctrl_retaddr(
	.clk(clk_clk),
	.d(\D_ctrl_retaddr~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_retaddr~q ),
	.prn(vcc));
defparam R_ctrl_retaddr.is_wysiwyg = "true";
defparam R_ctrl_retaddr.power_up = "low";

cyclone10lp_lcell_comb \R_src1~35 (
	.dataa(\R_ctrl_br~q ),
	.datab(\R_valid~q ),
	.datac(\R_ctrl_retaddr~q ),
	.datad(\E_valid_from_R~q ),
	.cin(gnd),
	.combout(\R_src1~35_combout ),
	.cout());
defparam \R_src1~35 .lut_mask = 16'hFFFE;
defparam \R_src1~35 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_src1[0]~37 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[0] ),
	.datad(\R_src1~35_combout ),
	.cin(gnd),
	.combout(\R_src1[0]~37_combout ),
	.cout());
defparam \R_src1[0]~37 .lut_mask = 16'hF7FF;
defparam \R_src1[0]~37 .sum_lutc_input = "datac";

dffeas \E_src1[0] (
	.clk(clk_clk),
	.d(\R_src1[0]~37_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[0]~q ),
	.prn(vcc));
defparam \E_src1[0] .is_wysiwyg = "true";
defparam \E_src1[0] .power_up = "low";

cyclone10lp_lcell_comb \Equal135~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\D_iw[10]~q ),
	.datad(\D_iw[9]~q ),
	.cin(gnd),
	.combout(\Equal135~0_combout ),
	.cout());
defparam \Equal135~0 .lut_mask = 16'h0FFF;
defparam \Equal135~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal135~1 (
	.dataa(\D_iw[7]~q ),
	.datab(\D_iw[6]~q ),
	.datac(\Equal135~0_combout ),
	.datad(\D_iw[8]~q ),
	.cin(gnd),
	.combout(\Equal135~1_combout ),
	.cout());
defparam \Equal135~1 .lut_mask = 16'hFEFF;
defparam \Equal135~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb D_op_wrctl(
	.dataa(\Equal0~9_combout ),
	.datab(\D_iw[14]~q ),
	.datac(\Equal62~13_combout ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_op_wrctl~combout ),
	.cout());
defparam D_op_wrctl.lut_mask = 16'hFEFF;
defparam D_op_wrctl.sum_lutc_input = "datac";

dffeas R_ctrl_wrctl_inst(
	.clk(clk_clk),
	.d(\D_op_wrctl~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_wrctl_inst~q ),
	.prn(vcc));
defparam R_ctrl_wrctl_inst.is_wysiwyg = "true";
defparam R_ctrl_wrctl_inst.power_up = "low";

cyclone10lp_lcell_comb \W_ienable_reg_nxt~0 (
	.dataa(\E_valid_from_R~q ),
	.datab(\Equal135~1_combout ),
	.datac(\R_ctrl_wrctl_inst~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\W_ienable_reg_nxt~0_combout ),
	.cout());
defparam \W_ienable_reg_nxt~0 .lut_mask = 16'hFEFE;
defparam \W_ienable_reg_nxt~0 .sum_lutc_input = "datac";

dffeas \W_ienable_reg[0] (
	.clk(clk_clk),
	.d(\E_src1[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_ienable_reg_nxt~0_combout ),
	.q(\W_ienable_reg[0]~q ),
	.prn(vcc));
defparam \W_ienable_reg[0] .is_wysiwyg = "true";
defparam \W_ienable_reg[0] .power_up = "low";

cyclone10lp_lcell_comb \W_ipending_reg_nxt[0]~0 (
	.dataa(\W_ienable_reg[0]~q ),
	.datab(av_readdata_9),
	.datac(av_readdata_8),
	.datad(\the_processor_nios2_gen2_0_cpu_nios2_oci|the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[0]~q ),
	.cin(gnd),
	.combout(\W_ipending_reg_nxt[0]~0_combout ),
	.cout());
defparam \W_ipending_reg_nxt[0]~0 .lut_mask = 16'hFEFF;
defparam \W_ipending_reg_nxt[0]~0 .sum_lutc_input = "datac";

dffeas \W_ipending_reg[0] (
	.clk(clk_clk),
	.d(\W_ipending_reg_nxt[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_ipending_reg[0]~q ),
	.prn(vcc));
defparam \W_ipending_reg[0] .is_wysiwyg = "true";
defparam \W_ipending_reg[0] .power_up = "low";

cyclone10lp_lcell_comb \R_src1[1]~36 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[1] ),
	.datad(\R_src1~35_combout ),
	.cin(gnd),
	.combout(\R_src1[1]~36_combout ),
	.cout());
defparam \R_src1[1]~36 .lut_mask = 16'hF7FF;
defparam \R_src1[1]~36 .sum_lutc_input = "datac";

dffeas \E_src1[1] (
	.clk(clk_clk),
	.d(\R_src1[1]~36_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[1]~q ),
	.prn(vcc));
defparam \E_src1[1] .is_wysiwyg = "true";
defparam \E_src1[1] .power_up = "low";

dffeas \W_ienable_reg[1] (
	.clk(clk_clk),
	.d(\E_src1[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_ienable_reg_nxt~0_combout ),
	.q(\W_ienable_reg[1]~q ),
	.prn(vcc));
defparam \W_ienable_reg[1] .is_wysiwyg = "true";
defparam \W_ienable_reg[1] .power_up = "low";

cyclone10lp_lcell_comb \W_ipending_reg_nxt[1]~1 (
	.dataa(\W_ienable_reg[1]~q ),
	.datab(irq),
	.datac(gnd),
	.datad(\the_processor_nios2_gen2_0_cpu_nios2_oci|the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[1]~q ),
	.cin(gnd),
	.combout(\W_ipending_reg_nxt[1]~1_combout ),
	.cout());
defparam \W_ipending_reg_nxt[1]~1 .lut_mask = 16'hEEFF;
defparam \W_ipending_reg_nxt[1]~1 .sum_lutc_input = "datac";

dffeas \W_ipending_reg[1] (
	.clk(clk_clk),
	.d(\W_ipending_reg_nxt[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_ipending_reg[1]~q ),
	.prn(vcc));
defparam \W_ipending_reg[1] .is_wysiwyg = "true";
defparam \W_ipending_reg[1] .power_up = "low";

cyclone10lp_lcell_comb \E_wrctl_status~1 (
	.dataa(\R_ctrl_wrctl_inst~q ),
	.datab(\D_iw[10]~q ),
	.datac(\D_iw[8]~q ),
	.datad(\D_iw[9]~q ),
	.cin(gnd),
	.combout(\E_wrctl_status~1_combout ),
	.cout());
defparam \E_wrctl_status~1 .lut_mask = 16'hBFFF;
defparam \E_wrctl_status~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_wrctl_estatus~0 (
	.dataa(\D_iw[6]~q ),
	.datab(\E_wrctl_status~1_combout ),
	.datac(gnd),
	.datad(\D_iw[7]~q ),
	.cin(gnd),
	.combout(\E_wrctl_estatus~0_combout ),
	.cout());
defparam \E_wrctl_estatus~0 .lut_mask = 16'hEEFF;
defparam \E_wrctl_estatus~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_exception~0 (
	.dataa(\Equal62~5_combout ),
	.datab(\D_op_opx_rsv63~0_combout ),
	.datac(\Equal62~6_combout ),
	.datad(\D_ctrl_implicit_dst_eretaddr~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~0_combout ),
	.cout());
defparam \D_ctrl_exception~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_exception~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_exception~1 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[12]~q ),
	.datac(\D_iw[13]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_exception~1_combout ),
	.cout());
defparam \D_ctrl_exception~1 .lut_mask = 16'hFBFF;
defparam \D_ctrl_exception~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_exception~2 (
	.dataa(\D_iw[16]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_ctrl_exception~2_combout ),
	.cout());
defparam \D_ctrl_exception~2 .lut_mask = 16'hAAFF;
defparam \D_ctrl_exception~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_exception~3 (
	.dataa(\Equal0~9_combout ),
	.datab(\D_ctrl_exception~0_combout ),
	.datac(\D_ctrl_exception~1_combout ),
	.datad(\D_ctrl_exception~2_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~3_combout ),
	.cout());
defparam \D_ctrl_exception~3 .lut_mask = 16'hFFFE;
defparam \D_ctrl_exception~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_implicit_dst_eretaddr~1 (
	.dataa(\D_iw[5]~q ),
	.datab(\Equal0~12_combout ),
	.datac(\Equal0~13_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~1_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~1 .lut_mask = 16'hFEFF;
defparam \D_ctrl_implicit_dst_eretaddr~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_implicit_dst_eretaddr~2 (
	.dataa(\Equal0~5_combout ),
	.datab(\Equal0~4_combout ),
	.datac(\Equal0~11_combout ),
	.datad(\D_ctrl_implicit_dst_eretaddr~1_combout ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~2_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~2 .lut_mask = 16'hBFFF;
defparam \D_ctrl_implicit_dst_eretaddr~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_implicit_dst_eretaddr~4 (
	.dataa(\D_ctrl_implicit_dst_eretaddr~2_combout ),
	.datab(\D_ctrl_implicit_dst_eretaddr~3_combout ),
	.datac(\Equal0~12_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~4_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~4 .lut_mask = 16'hEFFF;
defparam \D_ctrl_implicit_dst_eretaddr~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_exception~16 (
	.dataa(\D_ctrl_exception~3_combout ),
	.datab(\D_ctrl_exception~8_combout ),
	.datac(\D_ctrl_exception~15_combout ),
	.datad(\D_ctrl_implicit_dst_eretaddr~4_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~16_combout ),
	.cout());
defparam \D_ctrl_exception~16 .lut_mask = 16'hBFFF;
defparam \D_ctrl_exception~16 .sum_lutc_input = "datac";

dffeas R_ctrl_exception(
	.clk(clk_clk),
	.d(\D_ctrl_exception~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_exception~q ),
	.prn(vcc));
defparam R_ctrl_exception.is_wysiwyg = "true";
defparam R_ctrl_exception.power_up = "low";

cyclone10lp_lcell_comb \W_estatus_reg_inst_nxt~0 (
	.dataa(\E_src1[0]~q ),
	.datab(\W_estatus_reg~q ),
	.datac(\E_wrctl_estatus~0_combout ),
	.datad(\R_ctrl_exception~q ),
	.cin(gnd),
	.combout(\W_estatus_reg_inst_nxt~0_combout ),
	.cout());
defparam \W_estatus_reg_inst_nxt~0 .lut_mask = 16'hACFF;
defparam \W_estatus_reg_inst_nxt~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_estatus_reg_inst_nxt~1 (
	.dataa(\W_estatus_reg_inst_nxt~0_combout ),
	.datab(\R_ctrl_exception~q ),
	.datac(\W_status_reg_pie~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\W_estatus_reg_inst_nxt~1_combout ),
	.cout());
defparam \W_estatus_reg_inst_nxt~1 .lut_mask = 16'hFEFE;
defparam \W_estatus_reg_inst_nxt~1 .sum_lutc_input = "datac";

dffeas W_estatus_reg(
	.clk(clk_clk),
	.d(\W_estatus_reg_inst_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\E_valid_from_R~q ),
	.q(\W_estatus_reg~q ),
	.prn(vcc));
defparam W_estatus_reg.is_wysiwyg = "true";
defparam W_estatus_reg.power_up = "low";

cyclone10lp_lcell_comb \E_wrctl_bstatus~0 (
	.dataa(\D_iw[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\D_iw[6]~q ),
	.cin(gnd),
	.combout(\E_wrctl_bstatus~0_combout ),
	.cout());
defparam \E_wrctl_bstatus~0 .lut_mask = 16'hAAFF;
defparam \E_wrctl_bstatus~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_bstatus_reg_inst_nxt~0 (
	.dataa(\E_src1[0]~q ),
	.datab(\W_bstatus_reg~q ),
	.datac(\E_wrctl_status~1_combout ),
	.datad(\E_wrctl_bstatus~0_combout ),
	.cin(gnd),
	.combout(\W_bstatus_reg_inst_nxt~0_combout ),
	.cout());
defparam \W_bstatus_reg_inst_nxt~0 .lut_mask = 16'hEFFE;
defparam \W_bstatus_reg_inst_nxt~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_break~0 (
	.dataa(\D_iw[13]~q ),
	.datab(\D_iw[16]~q ),
	.datac(\D_op_opx_rsv17~0_combout ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\D_ctrl_break~0_combout ),
	.cout());
defparam \D_ctrl_break~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_break~0 .sum_lutc_input = "datac";

dffeas R_ctrl_break(
	.clk(clk_clk),
	.d(\D_ctrl_break~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_break~q ),
	.prn(vcc));
defparam R_ctrl_break.is_wysiwyg = "true";
defparam R_ctrl_break.power_up = "low";

cyclone10lp_lcell_comb \W_bstatus_reg_inst_nxt~1 (
	.dataa(\W_status_reg_pie~q ),
	.datab(\W_bstatus_reg_inst_nxt~0_combout ),
	.datac(gnd),
	.datad(\R_ctrl_break~q ),
	.cin(gnd),
	.combout(\W_bstatus_reg_inst_nxt~1_combout ),
	.cout());
defparam \W_bstatus_reg_inst_nxt~1 .lut_mask = 16'hAACC;
defparam \W_bstatus_reg_inst_nxt~1 .sum_lutc_input = "datac";

dffeas W_bstatus_reg(
	.clk(clk_clk),
	.d(\W_bstatus_reg_inst_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\E_valid_from_R~q ),
	.q(\W_bstatus_reg~q ),
	.prn(vcc));
defparam W_bstatus_reg.is_wysiwyg = "true";
defparam W_bstatus_reg.power_up = "low";

cyclone10lp_lcell_comb \E_wrctl_status~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\D_iw[7]~q ),
	.datad(\D_iw[6]~q ),
	.cin(gnd),
	.combout(\E_wrctl_status~0_combout ),
	.cout());
defparam \E_wrctl_status~0 .lut_mask = 16'h0FFF;
defparam \E_wrctl_status~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_status_reg_pie_inst_nxt~0 (
	.dataa(\E_src1[0]~q ),
	.datab(\W_status_reg_pie~q ),
	.datac(\E_wrctl_status~0_combout ),
	.datad(\E_wrctl_status~1_combout ),
	.cin(gnd),
	.combout(\W_status_reg_pie_inst_nxt~0_combout ),
	.cout());
defparam \W_status_reg_pie_inst_nxt~0 .lut_mask = 16'hEFFE;
defparam \W_status_reg_pie_inst_nxt~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_status_reg_pie_inst_nxt~1 (
	.dataa(\W_bstatus_reg~q ),
	.datab(\W_status_reg_pie_inst_nxt~0_combout ),
	.datac(\D_op_cmpge~0_combout ),
	.datad(\Equal62~4_combout ),
	.cin(gnd),
	.combout(\W_status_reg_pie_inst_nxt~1_combout ),
	.cout());
defparam \W_status_reg_pie_inst_nxt~1 .lut_mask = 16'hEFFE;
defparam \W_status_reg_pie_inst_nxt~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb D_op_eret(
	.dataa(\Equal0~9_combout ),
	.datab(\Equal62~4_combout ),
	.datac(\D_iw[14]~q ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_op_eret~combout ),
	.cout());
defparam D_op_eret.lut_mask = 16'hEFFF;
defparam D_op_eret.sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_pc_sel_nxt.10~1 (
	.dataa(\R_ctrl_exception~q ),
	.datab(\R_ctrl_break~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\F_pc_sel_nxt.10~1_combout ),
	.cout());
defparam \F_pc_sel_nxt.10~1 .lut_mask = 16'hEEEE;
defparam \F_pc_sel_nxt.10~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_status_reg_pie_inst_nxt~2 (
	.dataa(\W_estatus_reg~q ),
	.datab(\W_status_reg_pie_inst_nxt~1_combout ),
	.datac(\D_op_eret~combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\W_status_reg_pie_inst_nxt~2_combout ),
	.cout());
defparam \W_status_reg_pie_inst_nxt~2 .lut_mask = 16'hACFF;
defparam \W_status_reg_pie_inst_nxt~2 .sum_lutc_input = "datac";

dffeas W_status_reg_pie(
	.clk(clk_clk),
	.d(\W_status_reg_pie_inst_nxt~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\E_valid_from_R~q ),
	.q(\W_status_reg_pie~q ),
	.prn(vcc));
defparam W_status_reg_pie.is_wysiwyg = "true";
defparam W_status_reg_pie.power_up = "low";

cyclone10lp_lcell_comb \D_iw[26]~0 (
	.dataa(gnd),
	.datab(\W_ipending_reg[0]~q ),
	.datac(\W_ipending_reg[1]~q ),
	.datad(\W_status_reg_pie~q ),
	.cin(gnd),
	.combout(\D_iw[26]~0_combout ),
	.cout());
defparam \D_iw[26]~0 .lut_mask = 16'h3FFF;
defparam \D_iw[26]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_iw[26]~1 (
	.dataa(\D_iw[26]~0_combout ),
	.datab(hbreak_enabled1),
	.datac(gnd),
	.datad(\hbreak_req~0_combout ),
	.cin(gnd),
	.combout(\D_iw[26]~1_combout ),
	.cout());
defparam \D_iw[26]~1 .lut_mask = 16'hEEFF;
defparam \D_iw[26]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[1]~15 (
	.dataa(src1_valid),
	.datab(av_readdata_pre_1),
	.datac(gnd),
	.datad(\D_iw[26]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[1]~15_combout ),
	.cout());
defparam \F_iw[1]~15 .lut_mask = 16'hEEFF;
defparam \F_iw[1]~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[1]~16 (
	.dataa(src1_valid1),
	.datab(src1_valid2),
	.datac(q_a_1),
	.datad(av_readdata_pre_11),
	.cin(gnd),
	.combout(\F_iw[1]~16_combout ),
	.cout());
defparam \F_iw[1]~16 .lut_mask = 16'hFFFE;
defparam \F_iw[1]~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[1]~17 (
	.dataa(src1_valid3),
	.datab(src1_valid4),
	.datac(av_readdata_pre_12),
	.datad(av_readdata_pre_13),
	.cin(gnd),
	.combout(\F_iw[1]~17_combout ),
	.cout());
defparam \F_iw[1]~17 .lut_mask = 16'hFFFE;
defparam \F_iw[1]~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[1]~18 (
	.dataa(src_payload),
	.datab(src_payload1),
	.datac(av_readdata_pre_14),
	.datad(av_readdata_pre_15),
	.cin(gnd),
	.combout(\F_iw[1]~18_combout ),
	.cout());
defparam \F_iw[1]~18 .lut_mask = 16'hFFFE;
defparam \F_iw[1]~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[1]~19 (
	.dataa(\F_iw[1]~15_combout ),
	.datab(\F_iw[1]~16_combout ),
	.datac(\F_iw[1]~17_combout ),
	.datad(\F_iw[1]~18_combout ),
	.cin(gnd),
	.combout(\F_iw[1]~19_combout ),
	.cout());
defparam \F_iw[1]~19 .lut_mask = 16'hFFFE;
defparam \F_iw[1]~19 .sum_lutc_input = "datac";

dffeas \D_iw[1] (
	.clk(clk_clk),
	.d(\F_iw[1]~19_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[1]~q ),
	.prn(vcc));
defparam \D_iw[1] .is_wysiwyg = "true";
defparam \D_iw[1] .power_up = "low";

cyclone10lp_lcell_comb \Equal0~4 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~4_combout ),
	.cout());
defparam \Equal0~4 .lut_mask = 16'hFBFF;
defparam \Equal0~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_op_cmpge~0 (
	.dataa(\Equal0~4_combout ),
	.datab(\Equal0~5_combout ),
	.datac(\D_iw[14]~q ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_op_cmpge~0_combout ),
	.cout());
defparam \D_op_cmpge~0 .lut_mask = 16'hFEFF;
defparam \D_op_cmpge~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal0~6 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~6_combout ),
	.cout());
defparam \Equal0~6 .lut_mask = 16'hFFBF;
defparam \Equal0~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_alu_subtract~2 (
	.dataa(\D_iw[4]~q ),
	.datab(\Equal0~6_combout ),
	.datac(\Equal0~7_combout ),
	.datad(\D_ctrl_alu_force_xor~14_combout ),
	.cin(gnd),
	.combout(\D_ctrl_alu_subtract~2_combout ),
	.cout());
defparam \D_ctrl_alu_subtract~2 .lut_mask = 16'h27FF;
defparam \D_ctrl_alu_subtract~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_alu_subtract~3 (
	.dataa(\D_op_cmpge~0_combout ),
	.datab(\Equal62~0_combout ),
	.datac(gnd),
	.datad(\D_ctrl_alu_subtract~2_combout ),
	.cin(gnd),
	.combout(\D_ctrl_alu_subtract~3_combout ),
	.cout());
defparam \D_ctrl_alu_subtract~3 .lut_mask = 16'hEEFF;
defparam \D_ctrl_alu_subtract~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_alu_subtract~4 (
	.dataa(\Equal62~2_combout ),
	.datab(\Equal62~0_combout ),
	.datac(\Equal62~1_combout ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_alu_subtract~4_combout ),
	.cout());
defparam \D_ctrl_alu_subtract~4 .lut_mask = 16'hFAFC;
defparam \D_ctrl_alu_subtract~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_alu_subtract~5 (
	.dataa(\D_iw[14]~q ),
	.datab(\D_iw[15]~q ),
	.datac(\Equal62~1_combout ),
	.datad(\D_ctrl_alu_subtract~4_combout ),
	.cin(gnd),
	.combout(\D_ctrl_alu_subtract~5_combout ),
	.cout());
defparam \D_ctrl_alu_subtract~5 .lut_mask = 16'hFFB8;
defparam \D_ctrl_alu_subtract~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_alu_sub~0 (
	.dataa(\R_valid~q ),
	.datab(\D_ctrl_alu_subtract~3_combout ),
	.datac(\Equal0~9_combout ),
	.datad(\D_ctrl_alu_subtract~5_combout ),
	.cin(gnd),
	.combout(\E_alu_sub~0_combout ),
	.cout());
defparam \E_alu_sub~0 .lut_mask = 16'hFFFE;
defparam \E_alu_sub~0 .sum_lutc_input = "datac";

dffeas E_alu_sub(
	.clk(clk_clk),
	.d(\E_alu_sub~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_alu_sub~q ),
	.prn(vcc));
defparam E_alu_sub.is_wysiwyg = "true";
defparam E_alu_sub.power_up = "low";

cyclone10lp_lcell_comb \E_src2[13]~15 (
	.dataa(\R_ctrl_src_imm5_shift_rot~q ),
	.datab(\R_ctrl_hi_imm16~q ),
	.datac(\R_ctrl_force_src2_zero~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\E_src2[13]~15_combout ),
	.cout());
defparam \E_src2[13]~15 .lut_mask = 16'hFEFE;
defparam \E_src2[13]~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_src2_lo[7]~0 (
	.dataa(\D_iw[13]~q ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[13]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[7]~0_combout ),
	.cout());
defparam \R_src2_lo[7]~0 .lut_mask = 16'hACFF;
defparam \R_src2_lo[7]~0 .sum_lutc_input = "datac";

dffeas \E_src2[7] (
	.clk(clk_clk),
	.d(\R_src2_lo[7]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[7]~q ),
	.prn(vcc));
defparam \E_src2[7] .is_wysiwyg = "true";
defparam \E_src2[7] .power_up = "low";

cyclone10lp_lcell_comb \Add1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[7]~q ),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout());
defparam \Add1~0 .lut_mask = 16'h0FF0;
defparam \Add1~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_src1~34 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_valid_from_R~q ),
	.datad(\R_ctrl_jmp_direct~q ),
	.cin(gnd),
	.combout(\R_src1~34_combout ),
	.cout());
defparam \R_src1~34 .lut_mask = 16'h0FFF;
defparam \R_src1~34 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_src1[7]~9 (
	.dataa(\D_iw[11]~q ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[7] ),
	.datac(gnd),
	.datad(\R_src1~34_combout ),
	.cin(gnd),
	.combout(\E_src1[7]~9_combout ),
	.cout());
defparam \E_src1[7]~9 .lut_mask = 16'hAACC;
defparam \E_src1[7]~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_pc_plus_one[0]~0 (
	.dataa(F_pc_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\F_pc_plus_one[0]~0_combout ),
	.cout(\F_pc_plus_one[0]~1 ));
defparam \F_pc_plus_one[0]~0 .lut_mask = 16'h55AA;
defparam \F_pc_plus_one[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_pc_plus_one[1]~2 (
	.dataa(F_pc_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[0]~1 ),
	.combout(\F_pc_plus_one[1]~2_combout ),
	.cout(\F_pc_plus_one[1]~3 ));
defparam \F_pc_plus_one[1]~2 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[1]~2 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \F_pc_plus_one[2]~4 (
	.dataa(F_pc_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[1]~3 ),
	.combout(\F_pc_plus_one[2]~4_combout ),
	.cout(\F_pc_plus_one[2]~5 ));
defparam \F_pc_plus_one[2]~4 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[2]~4 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \F_pc_plus_one[3]~6 (
	.dataa(F_pc_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[2]~5 ),
	.combout(\F_pc_plus_one[3]~6_combout ),
	.cout(\F_pc_plus_one[3]~7 ));
defparam \F_pc_plus_one[3]~6 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[3]~6 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \F_pc_plus_one[4]~8 (
	.dataa(F_pc_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[3]~7 ),
	.combout(\F_pc_plus_one[4]~8_combout ),
	.cout(\F_pc_plus_one[4]~9 ));
defparam \F_pc_plus_one[4]~8 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[4]~8 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \F_pc_plus_one[5]~10 (
	.dataa(F_pc_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[4]~9 ),
	.combout(\F_pc_plus_one[5]~10_combout ),
	.cout(\F_pc_plus_one[5]~11 ));
defparam \F_pc_plus_one[5]~10 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[5]~10 .sum_lutc_input = "cin";

dffeas \E_src1[7] (
	.clk(clk_clk),
	.d(\E_src1[7]~9_combout ),
	.asdata(\F_pc_plus_one[5]~10_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~35_combout ),
	.ena(vcc),
	.q(\E_src1[7]~q ),
	.prn(vcc));
defparam \E_src1[7] .is_wysiwyg = "true";
defparam \E_src1[7] .power_up = "low";

cyclone10lp_lcell_comb \R_src2_lo[6]~1 (
	.dataa(\D_iw[12]~q ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[13]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[6]~1_combout ),
	.cout());
defparam \R_src2_lo[6]~1 .lut_mask = 16'hACFF;
defparam \R_src2_lo[6]~1 .sum_lutc_input = "datac";

dffeas \E_src2[6] (
	.clk(clk_clk),
	.d(\R_src2_lo[6]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[6]~q ),
	.prn(vcc));
defparam \E_src2[6] .is_wysiwyg = "true";
defparam \E_src2[6] .power_up = "low";

cyclone10lp_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[6]~q ),
	.cin(gnd),
	.combout(\Add1~1_combout ),
	.cout());
defparam \Add1~1 .lut_mask = 16'h0FF0;
defparam \Add1~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_src1[6]~10 (
	.dataa(\D_iw[10]~q ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[6] ),
	.datac(gnd),
	.datad(\R_src1~34_combout ),
	.cin(gnd),
	.combout(\E_src1[6]~10_combout ),
	.cout());
defparam \E_src1[6]~10 .lut_mask = 16'hAACC;
defparam \E_src1[6]~10 .sum_lutc_input = "datac";

dffeas \E_src1[6] (
	.clk(clk_clk),
	.d(\E_src1[6]~10_combout ),
	.asdata(\F_pc_plus_one[4]~8_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~35_combout ),
	.ena(vcc),
	.q(\E_src1[6]~q ),
	.prn(vcc));
defparam \E_src1[6] .is_wysiwyg = "true";
defparam \E_src1[6] .power_up = "low";

cyclone10lp_lcell_comb \R_src2_lo[5]~2 (
	.dataa(\D_iw[11]~q ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[13]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[5]~2_combout ),
	.cout());
defparam \R_src2_lo[5]~2 .lut_mask = 16'hACFF;
defparam \R_src2_lo[5]~2 .sum_lutc_input = "datac";

dffeas \E_src2[5] (
	.clk(clk_clk),
	.d(\R_src2_lo[5]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[5]~q ),
	.prn(vcc));
defparam \E_src2[5] .is_wysiwyg = "true";
defparam \E_src2[5] .power_up = "low";

cyclone10lp_lcell_comb \Add1~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[5]~q ),
	.cin(gnd),
	.combout(\Add1~2_combout ),
	.cout());
defparam \Add1~2 .lut_mask = 16'h0FF0;
defparam \Add1~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_src1[5]~11 (
	.dataa(\D_iw[9]~q ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[5] ),
	.datac(gnd),
	.datad(\R_src1~34_combout ),
	.cin(gnd),
	.combout(\E_src1[5]~11_combout ),
	.cout());
defparam \E_src1[5]~11 .lut_mask = 16'hAACC;
defparam \E_src1[5]~11 .sum_lutc_input = "datac";

dffeas \E_src1[5] (
	.clk(clk_clk),
	.d(\E_src1[5]~11_combout ),
	.asdata(\F_pc_plus_one[3]~6_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~35_combout ),
	.ena(vcc),
	.q(\E_src1[5]~q ),
	.prn(vcc));
defparam \E_src1[5] .is_wysiwyg = "true";
defparam \E_src1[5] .power_up = "low";

cyclone10lp_lcell_comb \Add1~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_src2[4]~q ),
	.datad(\E_alu_sub~q ),
	.cin(gnd),
	.combout(\Add1~3_combout ),
	.cout());
defparam \Add1~3 .lut_mask = 16'h0FF0;
defparam \Add1~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_src1[4]~12 (
	.dataa(\D_iw[8]~q ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[4] ),
	.datac(gnd),
	.datad(\R_src1~34_combout ),
	.cin(gnd),
	.combout(\E_src1[4]~12_combout ),
	.cout());
defparam \E_src1[4]~12 .lut_mask = 16'hAACC;
defparam \E_src1[4]~12 .sum_lutc_input = "datac";

dffeas \E_src1[4] (
	.clk(clk_clk),
	.d(\E_src1[4]~12_combout ),
	.asdata(\F_pc_plus_one[2]~4_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~35_combout ),
	.ena(vcc),
	.q(\E_src1[4]~q ),
	.prn(vcc));
defparam \E_src1[4] .is_wysiwyg = "true";
defparam \E_src1[4] .power_up = "low";

cyclone10lp_lcell_comb \Add1~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[3]~q ),
	.cin(gnd),
	.combout(\Add1~4_combout ),
	.cout());
defparam \Add1~4 .lut_mask = 16'h0FF0;
defparam \Add1~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_src1[3]~14 (
	.dataa(\D_iw[7]~q ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[3] ),
	.datac(gnd),
	.datad(\R_src1~34_combout ),
	.cin(gnd),
	.combout(\E_src1[3]~14_combout ),
	.cout());
defparam \E_src1[3]~14 .lut_mask = 16'hAACC;
defparam \E_src1[3]~14 .sum_lutc_input = "datac";

dffeas \E_src1[3] (
	.clk(clk_clk),
	.d(\E_src1[3]~14_combout ),
	.asdata(\F_pc_plus_one[1]~2_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~35_combout ),
	.ena(vcc),
	.q(\E_src1[3]~q ),
	.prn(vcc));
defparam \E_src1[3] .is_wysiwyg = "true";
defparam \E_src1[3] .power_up = "low";

cyclone10lp_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[2]~q ),
	.cin(gnd),
	.combout(\Add1~5_combout ),
	.cout());
defparam \Add1~5 .lut_mask = 16'h0FF0;
defparam \Add1~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_src1[2]~13 (
	.dataa(\D_iw[6]~q ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[2] ),
	.datac(gnd),
	.datad(\R_src1~34_combout ),
	.cin(gnd),
	.combout(\E_src1[2]~13_combout ),
	.cout());
defparam \E_src1[2]~13 .lut_mask = 16'hAACC;
defparam \E_src1[2]~13 .sum_lutc_input = "datac";

dffeas \E_src1[2] (
	.clk(clk_clk),
	.d(\E_src1[2]~13_combout ),
	.asdata(\F_pc_plus_one[0]~0_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~35_combout ),
	.ena(vcc),
	.q(\E_src1[2]~q ),
	.prn(vcc));
defparam \E_src1[2] .is_wysiwyg = "true";
defparam \E_src1[2] .power_up = "low";

cyclone10lp_lcell_comb \Add1~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[1]~q ),
	.cin(gnd),
	.combout(\Add1~6_combout ),
	.cout());
defparam \Add1~6 .lut_mask = 16'h0FF0;
defparam \Add1~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Add1~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[0]~q ),
	.cin(gnd),
	.combout(\Add1~7_combout ),
	.cout());
defparam \Add1~7 .lut_mask = 16'h0FF0;
defparam \Add1~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Add1~9 (
	.dataa(\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\Add1~9_cout ));
defparam \Add1~9 .lut_mask = 16'h00AA;
defparam \Add1~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Add1~10 (
	.dataa(\Add1~7_combout ),
	.datab(\E_src1[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~9_cout ),
	.combout(\Add1~10_combout ),
	.cout(\Add1~11 ));
defparam \Add1~10 .lut_mask = 16'h967F;
defparam \Add1~10 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add1~12 (
	.dataa(\Add1~6_combout ),
	.datab(\E_src1[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~11 ),
	.combout(\Add1~12_combout ),
	.cout(\Add1~13 ));
defparam \Add1~12 .lut_mask = 16'h96EF;
defparam \Add1~12 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add1~14 (
	.dataa(\Add1~5_combout ),
	.datab(\E_src1[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~13 ),
	.combout(\Add1~14_combout ),
	.cout(\Add1~15 ));
defparam \Add1~14 .lut_mask = 16'h967F;
defparam \Add1~14 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add1~16 (
	.dataa(\Add1~4_combout ),
	.datab(\E_src1[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~15 ),
	.combout(\Add1~16_combout ),
	.cout(\Add1~17 ));
defparam \Add1~16 .lut_mask = 16'h96EF;
defparam \Add1~16 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add1~18 (
	.dataa(\Add1~3_combout ),
	.datab(\E_src1[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~17 ),
	.combout(\Add1~18_combout ),
	.cout(\Add1~19 ));
defparam \Add1~18 .lut_mask = 16'h967F;
defparam \Add1~18 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add1~20 (
	.dataa(\Add1~2_combout ),
	.datab(\E_src1[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~19 ),
	.combout(\Add1~20_combout ),
	.cout(\Add1~21 ));
defparam \Add1~20 .lut_mask = 16'h96EF;
defparam \Add1~20 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add1~22 (
	.dataa(\Add1~1_combout ),
	.datab(\E_src1[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~21 ),
	.combout(\Add1~22_combout ),
	.cout(\Add1~23 ));
defparam \Add1~22 .lut_mask = 16'h967F;
defparam \Add1~22 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add1~24 (
	.dataa(\Add1~0_combout ),
	.datab(\E_src1[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~23 ),
	.combout(\Add1~24_combout ),
	.cout(\Add1~25 ));
defparam \Add1~24 .lut_mask = 16'h96EF;
defparam \Add1~24 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \D_logic_op_raw[1]~0 (
	.dataa(\D_iw[4]~q ),
	.datab(\D_iw[15]~q ),
	.datac(\Equal0~4_combout ),
	.datad(\D_iw[5]~q ),
	.cin(gnd),
	.combout(\D_logic_op_raw[1]~0_combout ),
	.cout());
defparam \D_logic_op_raw[1]~0 .lut_mask = 16'hEFFF;
defparam \D_logic_op_raw[1]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_alu_force_xor~10 (
	.dataa(\D_op_cmpge~0_combout ),
	.datab(\Equal62~0_combout ),
	.datac(\D_ctrl_alu_force_xor~14_combout ),
	.datad(\Equal0~5_combout ),
	.cin(gnd),
	.combout(\D_ctrl_alu_force_xor~10_combout ),
	.cout());
defparam \D_ctrl_alu_force_xor~10 .lut_mask = 16'hFEFF;
defparam \D_ctrl_alu_force_xor~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_alu_force_xor~11 (
	.dataa(\Equal0~6_combout ),
	.datab(\D_iw[5]~q ),
	.datac(\Equal0~7_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_alu_force_xor~11_combout ),
	.cout());
defparam \D_ctrl_alu_force_xor~11 .lut_mask = 16'hFEFF;
defparam \D_ctrl_alu_force_xor~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_alu_force_xor~13 (
	.dataa(\D_iw[14]~q ),
	.datab(\D_iw[15]~q ),
	.datac(\Equal62~0_combout ),
	.datad(\Equal62~1_combout ),
	.cin(gnd),
	.combout(\D_ctrl_alu_force_xor~13_combout ),
	.cout());
defparam \D_ctrl_alu_force_xor~13 .lut_mask = 16'hFFB8;
defparam \D_ctrl_alu_force_xor~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_alu_force_xor~12 (
	.dataa(\D_ctrl_alu_force_xor~10_combout ),
	.datab(\D_ctrl_alu_force_xor~11_combout ),
	.datac(\Equal0~9_combout ),
	.datad(\D_ctrl_alu_force_xor~13_combout ),
	.cin(gnd),
	.combout(\D_ctrl_alu_force_xor~12_combout ),
	.cout());
defparam \D_ctrl_alu_force_xor~12 .lut_mask = 16'hFFFE;
defparam \D_ctrl_alu_force_xor~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_logic_op[1]~0 (
	.dataa(\D_logic_op_raw[1]~0_combout ),
	.datab(\D_ctrl_alu_force_xor~12_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_logic_op[1]~0_combout ),
	.cout());
defparam \D_logic_op[1]~0 .lut_mask = 16'hEEEE;
defparam \D_logic_op[1]~0 .sum_lutc_input = "datac";

dffeas \R_logic_op[1] (
	.clk(clk_clk),
	.d(\D_logic_op[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_logic_op[1]~q ),
	.prn(vcc));
defparam \R_logic_op[1] .is_wysiwyg = "true";
defparam \R_logic_op[1] .power_up = "low";

cyclone10lp_lcell_comb \D_logic_op[0]~1 (
	.dataa(\D_ctrl_alu_force_xor~12_combout ),
	.datab(\D_iw[14]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\Equal0~9_combout ),
	.cin(gnd),
	.combout(\D_logic_op[0]~1_combout ),
	.cout());
defparam \D_logic_op[0]~1 .lut_mask = 16'hFAFC;
defparam \D_logic_op[0]~1 .sum_lutc_input = "datac";

dffeas \R_logic_op[0] (
	.clk(clk_clk),
	.d(\D_logic_op[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_logic_op[0]~q ),
	.prn(vcc));
defparam \R_logic_op[0] .is_wysiwyg = "true";
defparam \R_logic_op[0] .power_up = "low";

cyclone10lp_lcell_comb \E_logic_result[7]~0 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[7]~q ),
	.datac(\E_src1[7]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[7]~0_combout ),
	.cout());
defparam \E_logic_result[7]~0 .lut_mask = 16'h6996;
defparam \E_logic_result[7]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal0~16 (
	.dataa(\D_iw[13]~q ),
	.datab(gnd),
	.datac(\D_iw[11]~q ),
	.datad(\D_iw[16]~q ),
	.cin(gnd),
	.combout(\Equal0~16_combout ),
	.cout());
defparam \Equal0~16 .lut_mask = 16'hAFFF;
defparam \Equal0~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal0~17 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~17_combout ),
	.cout());
defparam \Equal0~17 .lut_mask = 16'hFFF7;
defparam \Equal0~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_logic~0 (
	.dataa(gnd),
	.datab(\D_iw[4]~q ),
	.datac(\Equal0~13_combout ),
	.datad(\Equal0~17_combout ),
	.cin(gnd),
	.combout(\D_ctrl_logic~0_combout ),
	.cout());
defparam \D_ctrl_logic~0 .lut_mask = 16'h3FFF;
defparam \D_ctrl_logic~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb D_ctrl_logic(
	.dataa(\Equal0~9_combout ),
	.datab(\D_iw[12]~q ),
	.datac(\Equal0~16_combout ),
	.datad(\D_ctrl_logic~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_logic~combout ),
	.cout());
defparam D_ctrl_logic.lut_mask = 16'hFEFF;
defparam D_ctrl_logic.sum_lutc_input = "datac";

dffeas R_ctrl_logic(
	.clk(clk_clk),
	.d(\D_ctrl_logic~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_logic~q ),
	.prn(vcc));
defparam R_ctrl_logic.is_wysiwyg = "true";
defparam R_ctrl_logic.power_up = "low";

cyclone10lp_lcell_comb \W_alu_result[7]~9 (
	.dataa(\Add1~24_combout ),
	.datab(\E_logic_result[7]~0_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[7]~9_combout ),
	.cout());
defparam \W_alu_result[7]~9 .lut_mask = 16'hAACC;
defparam \W_alu_result[7]~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_shift_rot_right~0 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[12]~q ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[16]~q ),
	.cin(gnd),
	.combout(\D_ctrl_shift_rot_right~0_combout ),
	.cout());
defparam \D_ctrl_shift_rot_right~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_shift_rot_right~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_shift_rot_right~1 (
	.dataa(\Equal0~9_combout ),
	.datab(\D_iw[14]~q ),
	.datac(\D_ctrl_shift_rot_right~0_combout ),
	.datad(\D_iw[13]~q ),
	.cin(gnd),
	.combout(\D_ctrl_shift_rot_right~1_combout ),
	.cout());
defparam \D_ctrl_shift_rot_right~1 .lut_mask = 16'hFEFF;
defparam \D_ctrl_shift_rot_right~1 .sum_lutc_input = "datac";

dffeas R_ctrl_shift_rot_right(
	.clk(clk_clk),
	.d(\D_ctrl_shift_rot_right~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_shift_rot_right~q ),
	.prn(vcc));
defparam R_ctrl_shift_rot_right.is_wysiwyg = "true";
defparam R_ctrl_shift_rot_right.power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[6]~12 (
	.dataa(\E_shift_rot_result[7]~q ),
	.datab(\E_shift_rot_result[5]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[6]~12_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[6]~12 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[6]~12 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[6] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[6]~12_combout ),
	.asdata(\E_src1[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[6]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[6] .is_wysiwyg = "true";
defparam \E_shift_rot_result[6] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[5]~11 (
	.dataa(\E_shift_rot_result[6]~q ),
	.datab(\E_shift_rot_result[4]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[5]~11_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[5]~11 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[5]~11 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[5] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[5]~11_combout ),
	.asdata(\E_src1[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[5]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[5] .is_wysiwyg = "true";
defparam \E_shift_rot_result[5] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[4]~10 (
	.dataa(\E_shift_rot_result[5]~q ),
	.datab(\E_shift_rot_result[3]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[4]~10_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[4]~10 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[4]~10 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[4] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[4]~10_combout ),
	.asdata(\E_src1[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[4]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[4] .is_wysiwyg = "true";
defparam \E_shift_rot_result[4] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[3]~14 (
	.dataa(\E_shift_rot_result[4]~q ),
	.datab(\E_shift_rot_result[2]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[3]~14_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[3]~14 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[3]~14 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[3] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[3]~14_combout ),
	.asdata(\E_src1[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[3]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[3] .is_wysiwyg = "true";
defparam \E_shift_rot_result[3] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[2]~13 (
	.dataa(\E_shift_rot_result[3]~q ),
	.datab(\E_shift_rot_result[1]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[2]~13_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[2]~13 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[2]~13 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[2] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[2]~13_combout ),
	.asdata(\E_src1[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[2]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[2] .is_wysiwyg = "true";
defparam \E_shift_rot_result[2] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[1]~16 (
	.dataa(\E_shift_rot_result[2]~q ),
	.datab(\E_shift_rot_result[0]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[1]~16_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[1]~16 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[1]~16 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[1] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[1]~16_combout ),
	.asdata(\E_src1[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[1]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[1] .is_wysiwyg = "true";
defparam \E_shift_rot_result[1] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[0]~17 (
	.dataa(\E_shift_rot_result[1]~q ),
	.datab(\E_shift_rot_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[0]~17_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[0]~17 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[0]~17 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[0] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[0]~17_combout ),
	.asdata(\E_src1[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[0]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[0] .is_wysiwyg = "true";
defparam \E_shift_rot_result[0] .power_up = "low";

cyclone10lp_lcell_comb \R_ctrl_rot_right_nxt~0 (
	.dataa(\Equal0~9_combout ),
	.datab(\D_iw[14]~q ),
	.datac(\Equal62~14_combout ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\R_ctrl_rot_right_nxt~0_combout ),
	.cout());
defparam \R_ctrl_rot_right_nxt~0 .lut_mask = 16'hFEFF;
defparam \R_ctrl_rot_right_nxt~0 .sum_lutc_input = "datac";

dffeas R_ctrl_rot_right(
	.clk(clk_clk),
	.d(\R_ctrl_rot_right_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_rot_right~q ),
	.prn(vcc));
defparam R_ctrl_rot_right.is_wysiwyg = "true";
defparam R_ctrl_rot_right.power_up = "low";

cyclone10lp_lcell_comb \D_ctrl_shift_logical~1 (
	.dataa(\D_ctrl_shift_logical~0_combout ),
	.datab(\D_iw[14]~q ),
	.datac(\Equal62~7_combout ),
	.datad(\Equal62~14_combout ),
	.cin(gnd),
	.combout(\D_ctrl_shift_logical~1_combout ),
	.cout());
defparam \D_ctrl_shift_logical~1 .lut_mask = 16'hFFB8;
defparam \D_ctrl_shift_logical~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_shift_logical~2 (
	.dataa(\Equal0~9_combout ),
	.datab(\D_iw[15]~q ),
	.datac(\D_ctrl_shift_logical~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_shift_logical~2_combout ),
	.cout());
defparam \D_ctrl_shift_logical~2 .lut_mask = 16'hFEFE;
defparam \D_ctrl_shift_logical~2 .sum_lutc_input = "datac";

dffeas R_ctrl_shift_logical(
	.clk(clk_clk),
	.d(\D_ctrl_shift_logical~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_shift_logical~q ),
	.prn(vcc));
defparam R_ctrl_shift_logical.is_wysiwyg = "true";
defparam R_ctrl_shift_logical.power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_fill_bit~0 (
	.dataa(\E_shift_rot_result[0]~q ),
	.datab(\E_shift_rot_result[31]~q ),
	.datac(\R_ctrl_rot_right~q ),
	.datad(\R_ctrl_shift_logical~q ),
	.cin(gnd),
	.combout(\E_shift_rot_fill_bit~0_combout ),
	.cout());
defparam \E_shift_rot_fill_bit~0 .lut_mask = 16'hACFF;
defparam \E_shift_rot_fill_bit~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[31]~19 (
	.dataa(\E_shift_rot_fill_bit~0_combout ),
	.datab(\E_shift_rot_result[30]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[31]~19_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[31]~19 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[31]~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_src1[31]~38 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[31] ),
	.datad(\R_src1~35_combout ),
	.cin(gnd),
	.combout(\R_src1[31]~38_combout ),
	.cout());
defparam \R_src1[31]~38 .lut_mask = 16'hF7FF;
defparam \R_src1[31]~38 .sum_lutc_input = "datac";

dffeas \E_src1[31] (
	.clk(clk_clk),
	.d(\R_src1[31]~38_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[31]~q ),
	.prn(vcc));
defparam \E_src1[31] .is_wysiwyg = "true";
defparam \E_src1[31] .power_up = "low";

dffeas \E_shift_rot_result[31] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[31]~19_combout ),
	.asdata(\E_src1[31]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[31]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[31] .is_wysiwyg = "true";
defparam \E_shift_rot_result[31] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[30]~21 (
	.dataa(\E_shift_rot_result[31]~q ),
	.datab(\E_shift_rot_result[29]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[30]~21_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[30]~21 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[30]~21 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_src1[30]~39 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[30] ),
	.datad(\R_src1~35_combout ),
	.cin(gnd),
	.combout(\R_src1[30]~39_combout ),
	.cout());
defparam \R_src1[30]~39 .lut_mask = 16'hF7FF;
defparam \R_src1[30]~39 .sum_lutc_input = "datac";

dffeas \E_src1[30] (
	.clk(clk_clk),
	.d(\R_src1[30]~39_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[30]~q ),
	.prn(vcc));
defparam \E_src1[30] .is_wysiwyg = "true";
defparam \E_src1[30] .power_up = "low";

dffeas \E_shift_rot_result[30] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[30]~21_combout ),
	.asdata(\E_src1[30]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[30]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[30] .is_wysiwyg = "true";
defparam \E_shift_rot_result[30] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[29]~22 (
	.dataa(\E_shift_rot_result[30]~q ),
	.datab(\E_shift_rot_result[28]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[29]~22_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[29]~22 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[29]~22 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_src1[29]~40 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[29] ),
	.datad(\R_src1~35_combout ),
	.cin(gnd),
	.combout(\R_src1[29]~40_combout ),
	.cout());
defparam \R_src1[29]~40 .lut_mask = 16'hF7FF;
defparam \R_src1[29]~40 .sum_lutc_input = "datac";

dffeas \E_src1[29] (
	.clk(clk_clk),
	.d(\R_src1[29]~40_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[29]~q ),
	.prn(vcc));
defparam \E_src1[29] .is_wysiwyg = "true";
defparam \E_src1[29] .power_up = "low";

dffeas \E_shift_rot_result[29] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[29]~22_combout ),
	.asdata(\E_src1[29]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[29]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[29] .is_wysiwyg = "true";
defparam \E_shift_rot_result[29] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[28]~23 (
	.dataa(\E_shift_rot_result[29]~q ),
	.datab(\E_shift_rot_result[27]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[28]~23_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[28]~23 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[28]~23 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_src1[28]~41 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[28] ),
	.datad(\R_src1~35_combout ),
	.cin(gnd),
	.combout(\R_src1[28]~41_combout ),
	.cout());
defparam \R_src1[28]~41 .lut_mask = 16'hF7FF;
defparam \R_src1[28]~41 .sum_lutc_input = "datac";

dffeas \E_src1[28] (
	.clk(clk_clk),
	.d(\R_src1[28]~41_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[28]~q ),
	.prn(vcc));
defparam \E_src1[28] .is_wysiwyg = "true";
defparam \E_src1[28] .power_up = "low";

dffeas \E_shift_rot_result[28] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[28]~23_combout ),
	.asdata(\E_src1[28]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[28]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[28] .is_wysiwyg = "true";
defparam \E_shift_rot_result[28] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[27]~24 (
	.dataa(\E_shift_rot_result[28]~q ),
	.datab(\E_shift_rot_result[26]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[27]~24_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[27]~24 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[27]~24 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_src1[27]~42 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[27] ),
	.datad(\R_src1~35_combout ),
	.cin(gnd),
	.combout(\R_src1[27]~42_combout ),
	.cout());
defparam \R_src1[27]~42 .lut_mask = 16'hF7FF;
defparam \R_src1[27]~42 .sum_lutc_input = "datac";

dffeas \E_src1[27] (
	.clk(clk_clk),
	.d(\R_src1[27]~42_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[27]~q ),
	.prn(vcc));
defparam \E_src1[27] .is_wysiwyg = "true";
defparam \E_src1[27] .power_up = "low";

dffeas \E_shift_rot_result[27] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[27]~24_combout ),
	.asdata(\E_src1[27]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[27]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[27] .is_wysiwyg = "true";
defparam \E_shift_rot_result[27] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[26]~25 (
	.dataa(\E_shift_rot_result[27]~q ),
	.datab(\E_shift_rot_result[25]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[26]~25_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[26]~25 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[26]~25 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_src1[26]~43 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[26] ),
	.datad(\R_src1~35_combout ),
	.cin(gnd),
	.combout(\R_src1[26]~43_combout ),
	.cout());
defparam \R_src1[26]~43 .lut_mask = 16'hF7FF;
defparam \R_src1[26]~43 .sum_lutc_input = "datac";

dffeas \E_src1[26] (
	.clk(clk_clk),
	.d(\R_src1[26]~43_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[26]~q ),
	.prn(vcc));
defparam \E_src1[26] .is_wysiwyg = "true";
defparam \E_src1[26] .power_up = "low";

dffeas \E_shift_rot_result[26] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[26]~25_combout ),
	.asdata(\E_src1[26]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[26]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[26] .is_wysiwyg = "true";
defparam \E_shift_rot_result[26] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[25]~26 (
	.dataa(\E_shift_rot_result[26]~q ),
	.datab(\E_shift_rot_result[24]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[25]~26_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[25]~26 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[25]~26 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_src1[25]~44 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[25] ),
	.datad(\R_src1~35_combout ),
	.cin(gnd),
	.combout(\R_src1[25]~44_combout ),
	.cout());
defparam \R_src1[25]~44 .lut_mask = 16'hF7FF;
defparam \R_src1[25]~44 .sum_lutc_input = "datac";

dffeas \E_src1[25] (
	.clk(clk_clk),
	.d(\R_src1[25]~44_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[25]~q ),
	.prn(vcc));
defparam \E_src1[25] .is_wysiwyg = "true";
defparam \E_src1[25] .power_up = "low";

dffeas \E_shift_rot_result[25] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[25]~26_combout ),
	.asdata(\E_src1[25]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[25]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[25] .is_wysiwyg = "true";
defparam \E_shift_rot_result[25] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[24]~27 (
	.dataa(\E_shift_rot_result[25]~q ),
	.datab(\E_shift_rot_result[23]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[24]~27_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[24]~27 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[24]~27 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_src1[24]~45 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[24] ),
	.datad(\R_src1~35_combout ),
	.cin(gnd),
	.combout(\R_src1[24]~45_combout ),
	.cout());
defparam \R_src1[24]~45 .lut_mask = 16'hF7FF;
defparam \R_src1[24]~45 .sum_lutc_input = "datac";

dffeas \E_src1[24] (
	.clk(clk_clk),
	.d(\R_src1[24]~45_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[24]~q ),
	.prn(vcc));
defparam \E_src1[24] .is_wysiwyg = "true";
defparam \E_src1[24] .power_up = "low";

dffeas \E_shift_rot_result[24] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[24]~27_combout ),
	.asdata(\E_src1[24]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[24]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[24] .is_wysiwyg = "true";
defparam \E_shift_rot_result[24] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[23]~28 (
	.dataa(\E_shift_rot_result[24]~q ),
	.datab(\E_shift_rot_result[22]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[23]~28_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[23]~28 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[23]~28 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_src1[23]~46 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[23] ),
	.datad(\R_src1~35_combout ),
	.cin(gnd),
	.combout(\R_src1[23]~46_combout ),
	.cout());
defparam \R_src1[23]~46 .lut_mask = 16'hF7FF;
defparam \R_src1[23]~46 .sum_lutc_input = "datac";

dffeas \E_src1[23] (
	.clk(clk_clk),
	.d(\R_src1[23]~46_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[23]~q ),
	.prn(vcc));
defparam \E_src1[23] .is_wysiwyg = "true";
defparam \E_src1[23] .power_up = "low";

dffeas \E_shift_rot_result[23] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[23]~28_combout ),
	.asdata(\E_src1[23]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[23]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[23] .is_wysiwyg = "true";
defparam \E_shift_rot_result[23] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[22]~29 (
	.dataa(\E_shift_rot_result[23]~q ),
	.datab(\E_shift_rot_result[21]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[22]~29_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[22]~29 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[22]~29 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_src1[22]~47 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[22] ),
	.datad(\R_src1~35_combout ),
	.cin(gnd),
	.combout(\R_src1[22]~47_combout ),
	.cout());
defparam \R_src1[22]~47 .lut_mask = 16'hF7FF;
defparam \R_src1[22]~47 .sum_lutc_input = "datac";

dffeas \E_src1[22] (
	.clk(clk_clk),
	.d(\R_src1[22]~47_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[22]~q ),
	.prn(vcc));
defparam \E_src1[22] .is_wysiwyg = "true";
defparam \E_src1[22] .power_up = "low";

dffeas \E_shift_rot_result[22] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[22]~29_combout ),
	.asdata(\E_src1[22]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[22]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[22] .is_wysiwyg = "true";
defparam \E_shift_rot_result[22] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[21]~30 (
	.dataa(\E_shift_rot_result[22]~q ),
	.datab(\E_shift_rot_result[20]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[21]~30_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[21]~30 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[21]~30 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_src1[21]~48 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[21] ),
	.datad(\R_src1~35_combout ),
	.cin(gnd),
	.combout(\R_src1[21]~48_combout ),
	.cout());
defparam \R_src1[21]~48 .lut_mask = 16'hF7FF;
defparam \R_src1[21]~48 .sum_lutc_input = "datac";

dffeas \E_src1[21] (
	.clk(clk_clk),
	.d(\R_src1[21]~48_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[21]~q ),
	.prn(vcc));
defparam \E_src1[21] .is_wysiwyg = "true";
defparam \E_src1[21] .power_up = "low";

dffeas \E_shift_rot_result[21] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[21]~30_combout ),
	.asdata(\E_src1[21]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[21]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[21] .is_wysiwyg = "true";
defparam \E_shift_rot_result[21] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[20]~31 (
	.dataa(\E_shift_rot_result[21]~q ),
	.datab(\E_shift_rot_result[19]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[20]~31_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[20]~31 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[20]~31 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_src1[20]~49 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[20] ),
	.datad(\R_src1~35_combout ),
	.cin(gnd),
	.combout(\R_src1[20]~49_combout ),
	.cout());
defparam \R_src1[20]~49 .lut_mask = 16'hF7FF;
defparam \R_src1[20]~49 .sum_lutc_input = "datac";

dffeas \E_src1[20] (
	.clk(clk_clk),
	.d(\R_src1[20]~49_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[20]~q ),
	.prn(vcc));
defparam \E_src1[20] .is_wysiwyg = "true";
defparam \E_src1[20] .power_up = "low";

dffeas \E_shift_rot_result[20] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[20]~31_combout ),
	.asdata(\E_src1[20]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[20]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[20] .is_wysiwyg = "true";
defparam \E_shift_rot_result[20] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[19]~20 (
	.dataa(\E_shift_rot_result[20]~q ),
	.datab(\E_shift_rot_result[18]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[19]~20_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[19]~20 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[19]~20 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_src1[19]~50 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[19] ),
	.datad(\R_src1~35_combout ),
	.cin(gnd),
	.combout(\R_src1[19]~50_combout ),
	.cout());
defparam \R_src1[19]~50 .lut_mask = 16'hF7FF;
defparam \R_src1[19]~50 .sum_lutc_input = "datac";

dffeas \E_src1[19] (
	.clk(clk_clk),
	.d(\R_src1[19]~50_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[19]~q ),
	.prn(vcc));
defparam \E_src1[19] .is_wysiwyg = "true";
defparam \E_src1[19] .power_up = "low";

dffeas \E_shift_rot_result[19] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[19]~20_combout ),
	.asdata(\E_src1[19]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[19]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[19] .is_wysiwyg = "true";
defparam \E_shift_rot_result[19] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[18]~18 (
	.dataa(\E_shift_rot_result[19]~q ),
	.datab(\E_shift_rot_result[17]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[18]~18_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[18]~18 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[18]~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_src1[18]~51 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[18] ),
	.datad(\R_src1~35_combout ),
	.cin(gnd),
	.combout(\R_src1[18]~51_combout ),
	.cout());
defparam \R_src1[18]~51 .lut_mask = 16'hF7FF;
defparam \R_src1[18]~51 .sum_lutc_input = "datac";

dffeas \E_src1[18] (
	.clk(clk_clk),
	.d(\R_src1[18]~51_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[18]~q ),
	.prn(vcc));
defparam \E_src1[18] .is_wysiwyg = "true";
defparam \E_src1[18] .power_up = "low";

dffeas \E_shift_rot_result[18] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[18]~18_combout ),
	.asdata(\E_src1[18]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[18]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[18] .is_wysiwyg = "true";
defparam \E_shift_rot_result[18] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[17]~15 (
	.dataa(\E_shift_rot_result[18]~q ),
	.datab(\E_shift_rot_result[16]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[17]~15_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[17]~15 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[17]~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_src1[17]~52 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[17] ),
	.datad(\R_src1~35_combout ),
	.cin(gnd),
	.combout(\R_src1[17]~52_combout ),
	.cout());
defparam \R_src1[17]~52 .lut_mask = 16'hF7FF;
defparam \R_src1[17]~52 .sum_lutc_input = "datac";

dffeas \E_src1[17] (
	.clk(clk_clk),
	.d(\R_src1[17]~52_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[17]~q ),
	.prn(vcc));
defparam \E_src1[17] .is_wysiwyg = "true";
defparam \E_src1[17] .power_up = "low";

dffeas \E_shift_rot_result[17] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[17]~15_combout ),
	.asdata(\E_src1[17]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[17]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[17] .is_wysiwyg = "true";
defparam \E_shift_rot_result[17] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[16]~1 (
	.dataa(\E_shift_rot_result[17]~q ),
	.datab(\E_shift_rot_result[15]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[16]~1_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[16]~1 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[16]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[20]~64 (
	.dataa(src1_valid1),
	.datab(src1_valid2),
	.datac(q_a_20),
	.datad(av_readdata_pre_201),
	.cin(gnd),
	.combout(\F_iw[20]~64_combout ),
	.cout());
defparam \F_iw[20]~64 .lut_mask = 16'hFFFE;
defparam \F_iw[20]~64 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[20]~65 (
	.dataa(\F_iw[20]~64_combout ),
	.datab(src1_valid),
	.datac(av_readdata_pre_20),
	.datad(\D_iw[26]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[20]~65_combout ),
	.cout());
defparam \F_iw[20]~65 .lut_mask = 16'hFEFF;
defparam \F_iw[20]~65 .sum_lutc_input = "datac";

dffeas \D_iw[20] (
	.clk(clk_clk),
	.d(\F_iw[20]~65_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[20]~q ),
	.prn(vcc));
defparam \D_iw[20] .is_wysiwyg = "true";
defparam \D_iw[20] .power_up = "low";

cyclone10lp_lcell_comb \E_src1[16]~0 (
	.dataa(\D_iw[20]~q ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[16] ),
	.datac(gnd),
	.datad(\R_src1~34_combout ),
	.cin(gnd),
	.combout(\E_src1[16]~0_combout ),
	.cout());
defparam \E_src1[16]~0 .lut_mask = 16'hAACC;
defparam \E_src1[16]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_pc_plus_one[6]~12 (
	.dataa(F_pc_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[5]~11 ),
	.combout(\F_pc_plus_one[6]~12_combout ),
	.cout(\F_pc_plus_one[6]~13 ));
defparam \F_pc_plus_one[6]~12 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[6]~12 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \F_pc_plus_one[7]~14 (
	.dataa(F_pc_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[6]~13 ),
	.combout(\F_pc_plus_one[7]~14_combout ),
	.cout(\F_pc_plus_one[7]~15 ));
defparam \F_pc_plus_one[7]~14 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[7]~14 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \F_pc_plus_one[8]~16 (
	.dataa(F_pc_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[7]~15 ),
	.combout(\F_pc_plus_one[8]~16_combout ),
	.cout(\F_pc_plus_one[8]~17 ));
defparam \F_pc_plus_one[8]~16 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[8]~16 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \F_pc_plus_one[9]~18 (
	.dataa(F_pc_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[8]~17 ),
	.combout(\F_pc_plus_one[9]~18_combout ),
	.cout(\F_pc_plus_one[9]~19 ));
defparam \F_pc_plus_one[9]~18 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[9]~18 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \F_pc_plus_one[10]~20 (
	.dataa(F_pc_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[9]~19 ),
	.combout(\F_pc_plus_one[10]~20_combout ),
	.cout(\F_pc_plus_one[10]~21 ));
defparam \F_pc_plus_one[10]~20 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[10]~20 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \F_pc_plus_one[11]~22 (
	.dataa(F_pc_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[10]~21 ),
	.combout(\F_pc_plus_one[11]~22_combout ),
	.cout(\F_pc_plus_one[11]~23 ));
defparam \F_pc_plus_one[11]~22 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[11]~22 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \F_pc_plus_one[12]~24 (
	.dataa(F_pc_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[11]~23 ),
	.combout(\F_pc_plus_one[12]~24_combout ),
	.cout(\F_pc_plus_one[12]~25 ));
defparam \F_pc_plus_one[12]~24 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[12]~24 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \F_pc_plus_one[13]~26 (
	.dataa(F_pc_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[12]~25 ),
	.combout(\F_pc_plus_one[13]~26_combout ),
	.cout(\F_pc_plus_one[13]~27 ));
defparam \F_pc_plus_one[13]~26 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[13]~26 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \F_pc_plus_one[14]~28 (
	.dataa(F_pc_14),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\F_pc_plus_one[13]~27 ),
	.combout(\F_pc_plus_one[14]~28_combout ),
	.cout());
defparam \F_pc_plus_one[14]~28 .lut_mask = 16'h5A5A;
defparam \F_pc_plus_one[14]~28 .sum_lutc_input = "cin";

dffeas \E_src1[16] (
	.clk(clk_clk),
	.d(\E_src1[16]~0_combout ),
	.asdata(\F_pc_plus_one[14]~28_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~35_combout ),
	.ena(vcc),
	.q(\E_src1[16]~q ),
	.prn(vcc));
defparam \E_src1[16] .is_wysiwyg = "true";
defparam \E_src1[16] .power_up = "low";

dffeas \E_shift_rot_result[16] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[16]~1_combout ),
	.asdata(\E_src1[16]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[16]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[16] .is_wysiwyg = "true";
defparam \E_shift_rot_result[16] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[15]~2 (
	.dataa(\E_shift_rot_result[16]~q ),
	.datab(\E_shift_rot_result[14]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[15]~2_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[15]~2 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[15]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[19]~66 (
	.dataa(src1_valid1),
	.datab(src1_valid2),
	.datac(q_a_19),
	.datad(av_readdata_pre_191),
	.cin(gnd),
	.combout(\F_iw[19]~66_combout ),
	.cout());
defparam \F_iw[19]~66 .lut_mask = 16'hFFFE;
defparam \F_iw[19]~66 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[19]~67 (
	.dataa(\F_iw[19]~66_combout ),
	.datab(src1_valid),
	.datac(av_readdata_pre_19),
	.datad(\D_iw[26]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[19]~67_combout ),
	.cout());
defparam \F_iw[19]~67 .lut_mask = 16'hFEFF;
defparam \F_iw[19]~67 .sum_lutc_input = "datac";

dffeas \D_iw[19] (
	.clk(clk_clk),
	.d(\F_iw[19]~67_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[19]~q ),
	.prn(vcc));
defparam \D_iw[19] .is_wysiwyg = "true";
defparam \D_iw[19] .power_up = "low";

cyclone10lp_lcell_comb \E_src1[15]~1 (
	.dataa(\D_iw[19]~q ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[15] ),
	.datac(gnd),
	.datad(\R_src1~34_combout ),
	.cin(gnd),
	.combout(\E_src1[15]~1_combout ),
	.cout());
defparam \E_src1[15]~1 .lut_mask = 16'hAACC;
defparam \E_src1[15]~1 .sum_lutc_input = "datac";

dffeas \E_src1[15] (
	.clk(clk_clk),
	.d(\E_src1[15]~1_combout ),
	.asdata(\F_pc_plus_one[13]~26_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~35_combout ),
	.ena(vcc),
	.q(\E_src1[15]~q ),
	.prn(vcc));
defparam \E_src1[15] .is_wysiwyg = "true";
defparam \E_src1[15] .power_up = "low";

dffeas \E_shift_rot_result[15] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[15]~2_combout ),
	.asdata(\E_src1[15]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[15]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[15] .is_wysiwyg = "true";
defparam \E_shift_rot_result[15] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[14]~3 (
	.dataa(\E_shift_rot_result[15]~q ),
	.datab(\E_shift_rot_result[13]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[14]~3_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[14]~3 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[14]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[18]~68 (
	.dataa(src1_valid),
	.datab(av_readdata_pre_18),
	.datac(src1_valid1),
	.datad(av_readdata_pre_181),
	.cin(gnd),
	.combout(\F_iw[18]~68_combout ),
	.cout());
defparam \F_iw[18]~68 .lut_mask = 16'hFFFE;
defparam \F_iw[18]~68 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[18]~69 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(src1_valid2),
	.datac(q_a_18),
	.datad(\F_iw[18]~68_combout ),
	.cin(gnd),
	.combout(\F_iw[18]~69_combout ),
	.cout());
defparam \F_iw[18]~69 .lut_mask = 16'hFFFE;
defparam \F_iw[18]~69 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[18]~70 (
	.dataa(\F_iw[18]~69_combout ),
	.datab(\hbreak_req~0_combout ),
	.datac(gnd),
	.datad(hbreak_enabled1),
	.cin(gnd),
	.combout(\F_iw[18]~70_combout ),
	.cout());
defparam \F_iw[18]~70 .lut_mask = 16'hEEFF;
defparam \F_iw[18]~70 .sum_lutc_input = "datac";

dffeas \D_iw[18] (
	.clk(clk_clk),
	.d(\F_iw[18]~70_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[18]~q ),
	.prn(vcc));
defparam \D_iw[18] .is_wysiwyg = "true";
defparam \D_iw[18] .power_up = "low";

cyclone10lp_lcell_comb \E_src1[14]~2 (
	.dataa(\D_iw[18]~q ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[14] ),
	.datac(gnd),
	.datad(\R_src1~34_combout ),
	.cin(gnd),
	.combout(\E_src1[14]~2_combout ),
	.cout());
defparam \E_src1[14]~2 .lut_mask = 16'hAACC;
defparam \E_src1[14]~2 .sum_lutc_input = "datac";

dffeas \E_src1[14] (
	.clk(clk_clk),
	.d(\E_src1[14]~2_combout ),
	.asdata(\F_pc_plus_one[12]~24_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~35_combout ),
	.ena(vcc),
	.q(\E_src1[14]~q ),
	.prn(vcc));
defparam \E_src1[14] .is_wysiwyg = "true";
defparam \E_src1[14] .power_up = "low";

dffeas \E_shift_rot_result[14] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[14]~3_combout ),
	.asdata(\E_src1[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[14]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[14] .is_wysiwyg = "true";
defparam \E_shift_rot_result[14] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[13]~4 (
	.dataa(\E_shift_rot_result[14]~q ),
	.datab(\E_shift_rot_result[12]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[13]~4_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[13]~4 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[13]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[17]~71 (
	.dataa(src1_valid),
	.datab(av_readdata_pre_17),
	.datac(src1_valid1),
	.datad(av_readdata_pre_171),
	.cin(gnd),
	.combout(\F_iw[17]~71_combout ),
	.cout());
defparam \F_iw[17]~71 .lut_mask = 16'hFFFE;
defparam \F_iw[17]~71 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[17]~72 (
	.dataa(src1_valid2),
	.datab(q_a_17),
	.datac(\F_iw[17]~71_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\F_iw[17]~72_combout ),
	.cout());
defparam \F_iw[17]~72 .lut_mask = 16'hFEFE;
defparam \F_iw[17]~72 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[17]~84 (
	.dataa(\D_iw[26]~0_combout ),
	.datab(hbreak_enabled1),
	.datac(\hbreak_req~0_combout ),
	.datad(\F_iw[17]~72_combout ),
	.cin(gnd),
	.combout(\F_iw[17]~84_combout ),
	.cout());
defparam \F_iw[17]~84 .lut_mask = 16'hFFDF;
defparam \F_iw[17]~84 .sum_lutc_input = "datac";

dffeas \D_iw[17] (
	.clk(clk_clk),
	.d(\F_iw[17]~84_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[17]~q ),
	.prn(vcc));
defparam \D_iw[17] .is_wysiwyg = "true";
defparam \D_iw[17] .power_up = "low";

cyclone10lp_lcell_comb \E_src1[13]~3 (
	.dataa(\D_iw[17]~q ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[13] ),
	.datac(gnd),
	.datad(\R_src1~34_combout ),
	.cin(gnd),
	.combout(\E_src1[13]~3_combout ),
	.cout());
defparam \E_src1[13]~3 .lut_mask = 16'hAACC;
defparam \E_src1[13]~3 .sum_lutc_input = "datac";

dffeas \E_src1[13] (
	.clk(clk_clk),
	.d(\E_src1[13]~3_combout ),
	.asdata(\F_pc_plus_one[11]~22_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~35_combout ),
	.ena(vcc),
	.q(\E_src1[13]~q ),
	.prn(vcc));
defparam \E_src1[13] .is_wysiwyg = "true";
defparam \E_src1[13] .power_up = "low";

dffeas \E_shift_rot_result[13] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[13]~4_combout ),
	.asdata(\E_src1[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[13]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[13] .is_wysiwyg = "true";
defparam \E_shift_rot_result[13] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[12]~5 (
	.dataa(\E_shift_rot_result[13]~q ),
	.datab(\E_shift_rot_result[11]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[12]~5_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[12]~5 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[12]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_src1[12]~4 (
	.dataa(\D_iw[16]~q ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[12] ),
	.datac(gnd),
	.datad(\R_src1~34_combout ),
	.cin(gnd),
	.combout(\E_src1[12]~4_combout ),
	.cout());
defparam \E_src1[12]~4 .lut_mask = 16'hAACC;
defparam \E_src1[12]~4 .sum_lutc_input = "datac";

dffeas \E_src1[12] (
	.clk(clk_clk),
	.d(\E_src1[12]~4_combout ),
	.asdata(\F_pc_plus_one[10]~20_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~35_combout ),
	.ena(vcc),
	.q(\E_src1[12]~q ),
	.prn(vcc));
defparam \E_src1[12] .is_wysiwyg = "true";
defparam \E_src1[12] .power_up = "low";

dffeas \E_shift_rot_result[12] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[12]~5_combout ),
	.asdata(\E_src1[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[12]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[12] .is_wysiwyg = "true";
defparam \E_shift_rot_result[12] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[11]~6 (
	.dataa(\E_shift_rot_result[12]~q ),
	.datab(\E_shift_rot_result[10]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[11]~6_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[11]~6 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[11]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_src1[11]~5 (
	.dataa(\D_iw[15]~q ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[11] ),
	.datac(gnd),
	.datad(\R_src1~34_combout ),
	.cin(gnd),
	.combout(\E_src1[11]~5_combout ),
	.cout());
defparam \E_src1[11]~5 .lut_mask = 16'hAACC;
defparam \E_src1[11]~5 .sum_lutc_input = "datac";

dffeas \E_src1[11] (
	.clk(clk_clk),
	.d(\E_src1[11]~5_combout ),
	.asdata(\F_pc_plus_one[9]~18_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~35_combout ),
	.ena(vcc),
	.q(\E_src1[11]~q ),
	.prn(vcc));
defparam \E_src1[11] .is_wysiwyg = "true";
defparam \E_src1[11] .power_up = "low";

dffeas \E_shift_rot_result[11] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[11]~6_combout ),
	.asdata(\E_src1[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[11]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[11] .is_wysiwyg = "true";
defparam \E_shift_rot_result[11] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[10]~7 (
	.dataa(\E_shift_rot_result[11]~q ),
	.datab(\E_shift_rot_result[9]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[10]~7_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[10]~7 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[10]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_src1[10]~6 (
	.dataa(\D_iw[14]~q ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[10] ),
	.datac(gnd),
	.datad(\R_src1~34_combout ),
	.cin(gnd),
	.combout(\E_src1[10]~6_combout ),
	.cout());
defparam \E_src1[10]~6 .lut_mask = 16'hAACC;
defparam \E_src1[10]~6 .sum_lutc_input = "datac";

dffeas \E_src1[10] (
	.clk(clk_clk),
	.d(\E_src1[10]~6_combout ),
	.asdata(\F_pc_plus_one[8]~16_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~35_combout ),
	.ena(vcc),
	.q(\E_src1[10]~q ),
	.prn(vcc));
defparam \E_src1[10] .is_wysiwyg = "true";
defparam \E_src1[10] .power_up = "low";

dffeas \E_shift_rot_result[10] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[10]~7_combout ),
	.asdata(\E_src1[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[10]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[10] .is_wysiwyg = "true";
defparam \E_shift_rot_result[10] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[9]~8 (
	.dataa(\E_shift_rot_result[10]~q ),
	.datab(\E_shift_rot_result[8]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[9]~8_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[9]~8 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[9]~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_src1[9]~7 (
	.dataa(\D_iw[13]~q ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[9] ),
	.datac(gnd),
	.datad(\R_src1~34_combout ),
	.cin(gnd),
	.combout(\E_src1[9]~7_combout ),
	.cout());
defparam \E_src1[9]~7 .lut_mask = 16'hAACC;
defparam \E_src1[9]~7 .sum_lutc_input = "datac";

dffeas \E_src1[9] (
	.clk(clk_clk),
	.d(\E_src1[9]~7_combout ),
	.asdata(\F_pc_plus_one[7]~14_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~35_combout ),
	.ena(vcc),
	.q(\E_src1[9]~q ),
	.prn(vcc));
defparam \E_src1[9] .is_wysiwyg = "true";
defparam \E_src1[9] .power_up = "low";

dffeas \E_shift_rot_result[9] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[9]~8_combout ),
	.asdata(\E_src1[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[9]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[9] .is_wysiwyg = "true";
defparam \E_shift_rot_result[9] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[8]~9 (
	.dataa(\E_shift_rot_result[9]~q ),
	.datab(\E_shift_rot_result[7]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[8]~9_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[8]~9 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[8]~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_src1[8]~8 (
	.dataa(\D_iw[12]~q ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[8] ),
	.datac(gnd),
	.datad(\R_src1~34_combout ),
	.cin(gnd),
	.combout(\E_src1[8]~8_combout ),
	.cout());
defparam \E_src1[8]~8 .lut_mask = 16'hAACC;
defparam \E_src1[8]~8 .sum_lutc_input = "datac";

dffeas \E_src1[8] (
	.clk(clk_clk),
	.d(\E_src1[8]~8_combout ),
	.asdata(\F_pc_plus_one[6]~12_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~35_combout ),
	.ena(vcc),
	.q(\E_src1[8]~q ),
	.prn(vcc));
defparam \E_src1[8] .is_wysiwyg = "true";
defparam \E_src1[8] .power_up = "low";

dffeas \E_shift_rot_result[8] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[8]~9_combout ),
	.asdata(\E_src1[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[8]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[8] .is_wysiwyg = "true";
defparam \E_shift_rot_result[8] .power_up = "low";

cyclone10lp_lcell_comb \E_shift_rot_result_nxt[7]~0 (
	.dataa(\E_shift_rot_result[8]~q ),
	.datab(\E_shift_rot_result[6]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[7]~0_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[7]~0 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[7]~0 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[7] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[7]~0_combout ),
	.asdata(\E_src1[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[7]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[7] .is_wysiwyg = "true";
defparam \E_shift_rot_result[7] .power_up = "low";

cyclone10lp_lcell_comb D_op_rdctl(
	.dataa(\Equal0~9_combout ),
	.datab(\Equal62~13_combout ),
	.datac(\D_iw[14]~q ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_op_rdctl~combout ),
	.cout());
defparam D_op_rdctl.lut_mask = 16'hEFFF;
defparam D_op_rdctl.sum_lutc_input = "datac";

dffeas R_ctrl_rd_ctl_reg(
	.clk(clk_clk),
	.d(\D_op_rdctl~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_rd_ctl_reg~q ),
	.prn(vcc));
defparam R_ctrl_rd_ctl_reg.is_wysiwyg = "true";
defparam R_ctrl_rd_ctl_reg.power_up = "low";

cyclone10lp_lcell_comb \Equal0~8 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~8_combout ),
	.cout());
defparam \Equal0~8 .lut_mask = 16'hF7FF;
defparam \Equal0~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_br_cmp~2 (
	.dataa(\Equal0~8_combout ),
	.datab(\Equal0~7_combout ),
	.datac(\Equal0~5_combout ),
	.datad(\D_ctrl_jmp_direct~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_br_cmp~2_combout ),
	.cout());
defparam \D_ctrl_br_cmp~2 .lut_mask = 16'hEFFF;
defparam \D_ctrl_br_cmp~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_br_cmp~5 (
	.dataa(\D_iw[14]~q ),
	.datab(\D_iw[15]~q ),
	.datac(\Equal62~0_combout ),
	.datad(\Equal62~1_combout ),
	.cin(gnd),
	.combout(\D_ctrl_br_cmp~5_combout ),
	.cout());
defparam \D_ctrl_br_cmp~5 .lut_mask = 16'hF7D5;
defparam \D_ctrl_br_cmp~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_br_cmp~3 (
	.dataa(\R_ctrl_br_nxt~1_combout ),
	.datab(\Equal0~9_combout ),
	.datac(\D_ctrl_br_cmp~5_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_br_cmp~3_combout ),
	.cout());
defparam \D_ctrl_br_cmp~3 .lut_mask = 16'hFEFE;
defparam \D_ctrl_br_cmp~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_br_cmp~4 (
	.dataa(\D_ctrl_br_cmp~2_combout ),
	.datab(\D_ctrl_br_cmp~3_combout ),
	.datac(\D_op_cmpge~0_combout ),
	.datad(\Equal62~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_br_cmp~4_combout ),
	.cout());
defparam \D_ctrl_br_cmp~4 .lut_mask = 16'hFFFE;
defparam \D_ctrl_br_cmp~4 .sum_lutc_input = "datac";

dffeas R_ctrl_br_cmp(
	.clk(clk_clk),
	.d(\D_ctrl_br_cmp~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_br_cmp~q ),
	.prn(vcc));
defparam R_ctrl_br_cmp.is_wysiwyg = "true";
defparam R_ctrl_br_cmp.power_up = "low";

cyclone10lp_lcell_comb \E_alu_result~0 (
	.dataa(\R_ctrl_rd_ctl_reg~q ),
	.datab(\R_ctrl_br_cmp~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\E_alu_result~0_combout ),
	.cout());
defparam \E_alu_result~0 .lut_mask = 16'hEEEE;
defparam \E_alu_result~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[21]~62 (
	.dataa(src1_valid1),
	.datab(src1_valid2),
	.datac(q_a_21),
	.datad(av_readdata_pre_211),
	.cin(gnd),
	.combout(\F_iw[21]~62_combout ),
	.cout());
defparam \F_iw[21]~62 .lut_mask = 16'hFFFE;
defparam \F_iw[21]~62 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_iw[21]~63 (
	.dataa(\F_iw[21]~62_combout ),
	.datab(src1_valid),
	.datac(av_readdata_pre_21),
	.datad(\D_iw[26]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[21]~63_combout ),
	.cout());
defparam \F_iw[21]~63 .lut_mask = 16'hFEFF;
defparam \F_iw[21]~63 .sum_lutc_input = "datac";

dffeas \D_iw[21] (
	.clk(clk_clk),
	.d(\F_iw[21]~63_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[21]~q ),
	.prn(vcc));
defparam \D_iw[21] .is_wysiwyg = "true";
defparam \D_iw[21] .power_up = "low";

cyclone10lp_lcell_comb \E_src2[16]~0 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[16]~0_combout ),
	.cout());
defparam \E_src2[16]~0 .lut_mask = 16'hAACC;
defparam \E_src2[16]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_unsigned_lo_imm16~3 (
	.dataa(\D_iw[5]~q ),
	.datab(\Equal0~7_combout ),
	.datac(\Equal0~8_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_unsigned_lo_imm16~3_combout ),
	.cout());
defparam \D_ctrl_unsigned_lo_imm16~3 .lut_mask = 16'hFAFC;
defparam \D_ctrl_unsigned_lo_imm16~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_unsigned_lo_imm16~4 (
	.dataa(\D_ctrl_unsigned_lo_imm16~5_combout ),
	.datab(\D_ctrl_unsigned_lo_imm16~3_combout ),
	.datac(\D_iw[5]~q ),
	.datad(\D_ctrl_logic~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_unsigned_lo_imm16~4_combout ),
	.cout());
defparam \D_ctrl_unsigned_lo_imm16~4 .lut_mask = 16'hEFFF;
defparam \D_ctrl_unsigned_lo_imm16~4 .sum_lutc_input = "datac";

dffeas R_ctrl_unsigned_lo_imm16(
	.clk(clk_clk),
	.d(\D_ctrl_unsigned_lo_imm16~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_unsigned_lo_imm16~q ),
	.prn(vcc));
defparam R_ctrl_unsigned_lo_imm16.is_wysiwyg = "true";
defparam R_ctrl_unsigned_lo_imm16.power_up = "low";

cyclone10lp_lcell_comb \R_src2_hi~0 (
	.dataa(\R_ctrl_force_src2_zero~q ),
	.datab(\R_ctrl_unsigned_lo_imm16~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\R_src2_hi~0_combout ),
	.cout());
defparam \R_src2_hi~0 .lut_mask = 16'hEEEE;
defparam \R_src2_hi~0 .sum_lutc_input = "datac";

dffeas \E_src2[16] (
	.clk(clk_clk),
	.d(\E_src2[16]~0_combout ),
	.asdata(\D_iw[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[16]~q ),
	.prn(vcc));
defparam \E_src2[16] .is_wysiwyg = "true";
defparam \E_src2[16] .power_up = "low";

cyclone10lp_lcell_comb \Add1~26 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[16]~q ),
	.cin(gnd),
	.combout(\Add1~26_combout ),
	.cout());
defparam \Add1~26 .lut_mask = 16'h0FF0;
defparam \Add1~26 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_src2_lo[15]~10 (
	.dataa(\D_iw[21]~q ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[13]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[15]~10_combout ),
	.cout());
defparam \R_src2_lo[15]~10 .lut_mask = 16'hACFF;
defparam \R_src2_lo[15]~10 .sum_lutc_input = "datac";

dffeas \E_src2[15] (
	.clk(clk_clk),
	.d(\R_src2_lo[15]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[15]~q ),
	.prn(vcc));
defparam \E_src2[15] .is_wysiwyg = "true";
defparam \E_src2[15] .power_up = "low";

cyclone10lp_lcell_comb \Add1~27 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[15]~q ),
	.cin(gnd),
	.combout(\Add1~27_combout ),
	.cout());
defparam \Add1~27 .lut_mask = 16'h0FF0;
defparam \Add1~27 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_src2_lo[14]~11 (
	.dataa(\D_iw[20]~q ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[13]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[14]~11_combout ),
	.cout());
defparam \R_src2_lo[14]~11 .lut_mask = 16'hACFF;
defparam \R_src2_lo[14]~11 .sum_lutc_input = "datac";

dffeas \E_src2[14] (
	.clk(clk_clk),
	.d(\R_src2_lo[14]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[14]~q ),
	.prn(vcc));
defparam \E_src2[14] .is_wysiwyg = "true";
defparam \E_src2[14] .power_up = "low";

cyclone10lp_lcell_comb \Add1~28 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[14]~q ),
	.cin(gnd),
	.combout(\Add1~28_combout ),
	.cout());
defparam \Add1~28 .lut_mask = 16'h0FF0;
defparam \Add1~28 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_src2_lo[13]~12 (
	.dataa(\D_iw[19]~q ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[13]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[13]~12_combout ),
	.cout());
defparam \R_src2_lo[13]~12 .lut_mask = 16'hACFF;
defparam \R_src2_lo[13]~12 .sum_lutc_input = "datac";

dffeas \E_src2[13] (
	.clk(clk_clk),
	.d(\R_src2_lo[13]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[13]~q ),
	.prn(vcc));
defparam \E_src2[13] .is_wysiwyg = "true";
defparam \E_src2[13] .power_up = "low";

cyclone10lp_lcell_comb \Add1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[13]~q ),
	.cin(gnd),
	.combout(\Add1~29_combout ),
	.cout());
defparam \Add1~29 .lut_mask = 16'h0FF0;
defparam \Add1~29 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_src2_lo[12]~13 (
	.dataa(\D_iw[18]~q ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[13]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[12]~13_combout ),
	.cout());
defparam \R_src2_lo[12]~13 .lut_mask = 16'hACFF;
defparam \R_src2_lo[12]~13 .sum_lutc_input = "datac";

dffeas \E_src2[12] (
	.clk(clk_clk),
	.d(\R_src2_lo[12]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[12]~q ),
	.prn(vcc));
defparam \E_src2[12] .is_wysiwyg = "true";
defparam \E_src2[12] .power_up = "low";

cyclone10lp_lcell_comb \Add1~30 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[12]~q ),
	.cin(gnd),
	.combout(\Add1~30_combout ),
	.cout());
defparam \Add1~30 .lut_mask = 16'h0FF0;
defparam \Add1~30 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_src2_lo[11]~14 (
	.dataa(\D_iw[17]~q ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[13]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[11]~14_combout ),
	.cout());
defparam \R_src2_lo[11]~14 .lut_mask = 16'hACFF;
defparam \R_src2_lo[11]~14 .sum_lutc_input = "datac";

dffeas \E_src2[11] (
	.clk(clk_clk),
	.d(\R_src2_lo[11]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[11]~q ),
	.prn(vcc));
defparam \E_src2[11] .is_wysiwyg = "true";
defparam \E_src2[11] .power_up = "low";

cyclone10lp_lcell_comb \Add1~31 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[11]~q ),
	.cin(gnd),
	.combout(\Add1~31_combout ),
	.cout());
defparam \Add1~31 .lut_mask = 16'h0FF0;
defparam \Add1~31 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_src2_lo[10]~15 (
	.dataa(\D_iw[16]~q ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[13]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[10]~15_combout ),
	.cout());
defparam \R_src2_lo[10]~15 .lut_mask = 16'hACFF;
defparam \R_src2_lo[10]~15 .sum_lutc_input = "datac";

dffeas \E_src2[10] (
	.clk(clk_clk),
	.d(\R_src2_lo[10]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[10]~q ),
	.prn(vcc));
defparam \E_src2[10] .is_wysiwyg = "true";
defparam \E_src2[10] .power_up = "low";

cyclone10lp_lcell_comb \Add1~32 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[10]~q ),
	.cin(gnd),
	.combout(\Add1~32_combout ),
	.cout());
defparam \Add1~32 .lut_mask = 16'h0FF0;
defparam \Add1~32 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_src2_lo[9]~16 (
	.dataa(\D_iw[15]~q ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[13]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[9]~16_combout ),
	.cout());
defparam \R_src2_lo[9]~16 .lut_mask = 16'hACFF;
defparam \R_src2_lo[9]~16 .sum_lutc_input = "datac";

dffeas \E_src2[9] (
	.clk(clk_clk),
	.d(\R_src2_lo[9]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[9]~q ),
	.prn(vcc));
defparam \E_src2[9] .is_wysiwyg = "true";
defparam \E_src2[9] .power_up = "low";

cyclone10lp_lcell_comb \Add1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[9]~q ),
	.cin(gnd),
	.combout(\Add1~33_combout ),
	.cout());
defparam \Add1~33 .lut_mask = 16'h0FF0;
defparam \Add1~33 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_src2_lo[8]~17 (
	.dataa(\D_iw[14]~q ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[13]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[8]~17_combout ),
	.cout());
defparam \R_src2_lo[8]~17 .lut_mask = 16'hACFF;
defparam \R_src2_lo[8]~17 .sum_lutc_input = "datac";

dffeas \E_src2[8] (
	.clk(clk_clk),
	.d(\R_src2_lo[8]~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[8]~q ),
	.prn(vcc));
defparam \E_src2[8] .is_wysiwyg = "true";
defparam \E_src2[8] .power_up = "low";

cyclone10lp_lcell_comb \Add1~34 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[8]~q ),
	.cin(gnd),
	.combout(\Add1~34_combout ),
	.cout());
defparam \Add1~34 .lut_mask = 16'h0FF0;
defparam \Add1~34 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Add1~35 (
	.dataa(\Add1~34_combout ),
	.datab(\E_src1[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~25 ),
	.combout(\Add1~35_combout ),
	.cout(\Add1~36 ));
defparam \Add1~35 .lut_mask = 16'h967F;
defparam \Add1~35 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add1~37 (
	.dataa(\Add1~33_combout ),
	.datab(\E_src1[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~36 ),
	.combout(\Add1~37_combout ),
	.cout(\Add1~38 ));
defparam \Add1~37 .lut_mask = 16'h96EF;
defparam \Add1~37 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add1~39 (
	.dataa(\Add1~32_combout ),
	.datab(\E_src1[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~38 ),
	.combout(\Add1~39_combout ),
	.cout(\Add1~40 ));
defparam \Add1~39 .lut_mask = 16'h967F;
defparam \Add1~39 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add1~41 (
	.dataa(\Add1~31_combout ),
	.datab(\E_src1[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~40 ),
	.combout(\Add1~41_combout ),
	.cout(\Add1~42 ));
defparam \Add1~41 .lut_mask = 16'h96EF;
defparam \Add1~41 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add1~43 (
	.dataa(\Add1~30_combout ),
	.datab(\E_src1[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~42 ),
	.combout(\Add1~43_combout ),
	.cout(\Add1~44 ));
defparam \Add1~43 .lut_mask = 16'h967F;
defparam \Add1~43 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add1~45 (
	.dataa(\Add1~29_combout ),
	.datab(\E_src1[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~44 ),
	.combout(\Add1~45_combout ),
	.cout(\Add1~46 ));
defparam \Add1~45 .lut_mask = 16'h96EF;
defparam \Add1~45 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add1~47 (
	.dataa(\Add1~28_combout ),
	.datab(\E_src1[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~46 ),
	.combout(\Add1~47_combout ),
	.cout(\Add1~48 ));
defparam \Add1~47 .lut_mask = 16'h967F;
defparam \Add1~47 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add1~49 (
	.dataa(\Add1~27_combout ),
	.datab(\E_src1[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~48 ),
	.combout(\Add1~49_combout ),
	.cout(\Add1~50 ));
defparam \Add1~49 .lut_mask = 16'h96EF;
defparam \Add1~49 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Add1~51 (
	.dataa(\Add1~26_combout ),
	.datab(\E_src1[16]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~50 ),
	.combout(\Add1~51_combout ),
	.cout(\Add1~52 ));
defparam \Add1~51 .lut_mask = 16'h967F;
defparam \Add1~51 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \E_logic_result[16]~1 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[16]~q ),
	.datac(\E_src1[16]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[16]~1_combout ),
	.cout());
defparam \E_logic_result[16]~1 .lut_mask = 16'h6996;
defparam \E_logic_result[16]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_alu_result[16]~0 (
	.dataa(\Add1~51_combout ),
	.datab(\E_logic_result[16]~1_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[16]~0_combout ),
	.cout());
defparam \W_alu_result[16]~0 .lut_mask = 16'hAACC;
defparam \W_alu_result[16]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_logic_result[15]~2 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[15]~q ),
	.datac(\E_src1[15]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[15]~2_combout ),
	.cout());
defparam \E_logic_result[15]~2 .lut_mask = 16'h6996;
defparam \E_logic_result[15]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_alu_result[15]~1 (
	.dataa(\Add1~49_combout ),
	.datab(\E_logic_result[15]~2_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[15]~1_combout ),
	.cout());
defparam \W_alu_result[15]~1 .lut_mask = 16'hAACC;
defparam \W_alu_result[15]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_logic_result[14]~3 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[14]~q ),
	.datac(\E_src1[14]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[14]~3_combout ),
	.cout());
defparam \E_logic_result[14]~3 .lut_mask = 16'h6996;
defparam \E_logic_result[14]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_alu_result[14]~2 (
	.dataa(\Add1~47_combout ),
	.datab(\E_logic_result[14]~3_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[14]~2_combout ),
	.cout());
defparam \W_alu_result[14]~2 .lut_mask = 16'hAACC;
defparam \W_alu_result[14]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_logic_result[13]~4 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[13]~q ),
	.datac(\E_src1[13]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[13]~4_combout ),
	.cout());
defparam \E_logic_result[13]~4 .lut_mask = 16'h6996;
defparam \E_logic_result[13]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_alu_result[13]~3 (
	.dataa(\Add1~45_combout ),
	.datab(\E_logic_result[13]~4_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[13]~3_combout ),
	.cout());
defparam \W_alu_result[13]~3 .lut_mask = 16'hAACC;
defparam \W_alu_result[13]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_logic_result[12]~5 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[12]~q ),
	.datac(\E_src1[12]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[12]~5_combout ),
	.cout());
defparam \E_logic_result[12]~5 .lut_mask = 16'h6996;
defparam \E_logic_result[12]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_alu_result[12]~4 (
	.dataa(\Add1~43_combout ),
	.datab(\E_logic_result[12]~5_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[12]~4_combout ),
	.cout());
defparam \W_alu_result[12]~4 .lut_mask = 16'hAACC;
defparam \W_alu_result[12]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_logic_result[11]~6 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[11]~q ),
	.datac(\E_src1[11]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[11]~6_combout ),
	.cout());
defparam \E_logic_result[11]~6 .lut_mask = 16'h6996;
defparam \E_logic_result[11]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_alu_result[11]~5 (
	.dataa(\Add1~41_combout ),
	.datab(\E_logic_result[11]~6_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[11]~5_combout ),
	.cout());
defparam \W_alu_result[11]~5 .lut_mask = 16'hAACC;
defparam \W_alu_result[11]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_logic_result[10]~7 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[10]~q ),
	.datac(\E_src1[10]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[10]~7_combout ),
	.cout());
defparam \E_logic_result[10]~7 .lut_mask = 16'h6996;
defparam \E_logic_result[10]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_alu_result[10]~6 (
	.dataa(\Add1~39_combout ),
	.datab(\E_logic_result[10]~7_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[10]~6_combout ),
	.cout());
defparam \W_alu_result[10]~6 .lut_mask = 16'hAACC;
defparam \W_alu_result[10]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_logic_result[9]~8 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[9]~q ),
	.datac(\E_src1[9]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[9]~8_combout ),
	.cout());
defparam \E_logic_result[9]~8 .lut_mask = 16'h6996;
defparam \E_logic_result[9]~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_alu_result[9]~7 (
	.dataa(\Add1~37_combout ),
	.datab(\E_logic_result[9]~8_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[9]~7_combout ),
	.cout());
defparam \W_alu_result[9]~7 .lut_mask = 16'hAACC;
defparam \W_alu_result[9]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_logic_result[8]~9 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[8]~q ),
	.datac(\E_src1[8]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[8]~9_combout ),
	.cout());
defparam \E_logic_result[8]~9 .lut_mask = 16'h6996;
defparam \E_logic_result[8]~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_alu_result[8]~8 (
	.dataa(\Add1~35_combout ),
	.datab(\E_logic_result[8]~9_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[8]~8_combout ),
	.cout());
defparam \W_alu_result[8]~8 .lut_mask = 16'hAACC;
defparam \W_alu_result[8]~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_logic_result[4]~10 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[4]~q ),
	.datac(\E_src1[4]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[4]~10_combout ),
	.cout());
defparam \E_logic_result[4]~10 .lut_mask = 16'h6996;
defparam \E_logic_result[4]~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_alu_result[4]~12 (
	.dataa(\Add1~18_combout ),
	.datab(\E_logic_result[4]~10_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[4]~12_combout ),
	.cout());
defparam \W_alu_result[4]~12 .lut_mask = 16'hAACC;
defparam \W_alu_result[4]~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_logic_result[5]~11 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[5]~q ),
	.datac(\E_src1[5]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[5]~11_combout ),
	.cout());
defparam \E_logic_result[5]~11 .lut_mask = 16'h6996;
defparam \E_logic_result[5]~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_alu_result[5]~11 (
	.dataa(\Add1~20_combout ),
	.datab(\E_logic_result[5]~11_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[5]~11_combout ),
	.cout());
defparam \W_alu_result[5]~11 .lut_mask = 16'hAACC;
defparam \W_alu_result[5]~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_logic_result[6]~12 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[6]~q ),
	.datac(\E_src1[6]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[6]~12_combout ),
	.cout());
defparam \E_logic_result[6]~12 .lut_mask = 16'h6996;
defparam \E_logic_result[6]~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_alu_result[6]~10 (
	.dataa(\Add1~22_combout ),
	.datab(\E_logic_result[6]~12_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[6]~10_combout ),
	.cout());
defparam \W_alu_result[6]~10 .lut_mask = 16'hAACC;
defparam \W_alu_result[6]~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_logic_result[2]~13 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[2]~q ),
	.datac(\E_src1[2]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[2]~13_combout ),
	.cout());
defparam \E_logic_result[2]~13 .lut_mask = 16'h6996;
defparam \E_logic_result[2]~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_alu_result[2]~13 (
	.dataa(\Add1~14_combout ),
	.datab(\E_logic_result[2]~13_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[2]~13_combout ),
	.cout());
defparam \W_alu_result[2]~13 .lut_mask = 16'hAACC;
defparam \W_alu_result[2]~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_logic_result[3]~14 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[3]~q ),
	.datac(\E_src1[3]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[3]~14_combout ),
	.cout());
defparam \E_logic_result[3]~14 .lut_mask = 16'h6996;
defparam \E_logic_result[3]~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \W_alu_result[3]~14 (
	.dataa(\Add1~16_combout ),
	.datab(\E_logic_result[3]~14_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[3]~14_combout ),
	.cout());
defparam \W_alu_result[3]~14 .lut_mask = 16'hAACC;
defparam \W_alu_result[3]~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_mem16~1 (
	.dataa(\D_ctrl_mem16~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_mem16~1_combout ),
	.cout());
defparam \D_ctrl_mem16~1 .lut_mask = 16'hAAFF;
defparam \D_ctrl_mem16~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \d_writedata[24]~0 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[24]~0_combout ),
	.cout());
defparam \d_writedata[24]~0 .lut_mask = 16'hAACC;
defparam \d_writedata[24]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_mem8~0 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[2]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_mem8~0_combout ),
	.cout());
defparam \D_ctrl_mem8~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_mem8~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_mem8~1 (
	.dataa(\D_ctrl_mem8~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_mem8~1_combout ),
	.cout());
defparam \D_ctrl_mem8~1 .lut_mask = 16'hAAFF;
defparam \D_ctrl_mem8~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \d_writedata[25]~1 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[25]~1_combout ),
	.cout());
defparam \d_writedata[25]~1 .lut_mask = 16'hAACC;
defparam \d_writedata[25]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \d_writedata[26]~2 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[26]~2_combout ),
	.cout());
defparam \d_writedata[26]~2 .lut_mask = 16'hAACC;
defparam \d_writedata[26]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \d_writedata[27]~3 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[27]~3_combout ),
	.cout());
defparam \d_writedata[27]~3 .lut_mask = 16'hAACC;
defparam \d_writedata[27]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \d_writedata[28]~4 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[28]~4_combout ),
	.cout());
defparam \d_writedata[28]~4 .lut_mask = 16'hAACC;
defparam \d_writedata[28]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \d_writedata[29]~5 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[29]~5_combout ),
	.cout());
defparam \d_writedata[29]~5 .lut_mask = 16'hAACC;
defparam \d_writedata[29]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \d_writedata[30]~6 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[30]~6_combout ),
	.cout());
defparam \d_writedata[30]~6 .lut_mask = 16'hAACC;
defparam \d_writedata[30]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \d_writedata[31]~7 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[31]~7_combout ),
	.cout());
defparam \d_writedata[31]~7 .lut_mask = 16'hAACC;
defparam \d_writedata[31]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \i_read_nxt~0 (
	.dataa(\W_valid~q ),
	.datab(i_read1),
	.datac(WideOr13),
	.datad(WideOr14),
	.cin(gnd),
	.combout(\i_read_nxt~0_combout ),
	.cout());
defparam \i_read_nxt~0 .lut_mask = 16'hFFFD;
defparam \i_read_nxt~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_uncond_cti_non_br~0 (
	.dataa(\Equal0~9_combout ),
	.datab(\Equal62~3_combout ),
	.datac(\D_iw[14]~q ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_ctrl_uncond_cti_non_br~0_combout ),
	.cout());
defparam \D_ctrl_uncond_cti_non_br~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_uncond_cti_non_br~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_ctrl_uncond_cti_non_br~2 (
	.dataa(\D_ctrl_jmp_direct~1_combout ),
	.datab(\D_ctrl_uncond_cti_non_br~0_combout ),
	.datac(gnd),
	.datad(\D_ctrl_uncond_cti_non_br~1_combout ),
	.cin(gnd),
	.combout(\D_ctrl_uncond_cti_non_br~2_combout ),
	.cout());
defparam \D_ctrl_uncond_cti_non_br~2 .lut_mask = 16'hEEFF;
defparam \D_ctrl_uncond_cti_non_br~2 .sum_lutc_input = "datac";

dffeas R_ctrl_uncond_cti_non_br(
	.clk(clk_clk),
	.d(\D_ctrl_uncond_cti_non_br~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_uncond_cti_non_br~q ),
	.prn(vcc));
defparam R_ctrl_uncond_cti_non_br.is_wysiwyg = "true";
defparam R_ctrl_uncond_cti_non_br.power_up = "low";

cyclone10lp_lcell_comb \Equal0~22 (
	.dataa(\D_iw[4]~q ),
	.datab(\D_iw[5]~q ),
	.datac(\Equal0~6_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal0~22_combout ),
	.cout());
defparam \Equal0~22 .lut_mask = 16'hF7F7;
defparam \Equal0~22 .sum_lutc_input = "datac";

dffeas R_ctrl_br_uncond(
	.clk(clk_clk),
	.d(\Equal0~22_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_br_uncond~q ),
	.prn(vcc));
defparam R_ctrl_br_uncond.is_wysiwyg = "true";
defparam R_ctrl_br_uncond.power_up = "low";

dffeas \R_compare_op[1] (
	.clk(clk_clk),
	.d(\D_logic_op_raw[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_compare_op[1]~q ),
	.prn(vcc));
defparam \R_compare_op[1] .is_wysiwyg = "true";
defparam \R_compare_op[1] .power_up = "low";

cyclone10lp_lcell_comb \R_src2_hi[15]~1 (
	.dataa(\D_iw[21]~q ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\R_ctrl_hi_imm16~q ),
	.cin(gnd),
	.combout(\R_src2_hi[15]~1_combout ),
	.cout());
defparam \R_src2_hi[15]~1 .lut_mask = 16'hEFFE;
defparam \R_src2_hi[15]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \R_src2_hi[15]~2 (
	.dataa(\R_src2_hi[15]~1_combout ),
	.datab(gnd),
	.datac(\R_ctrl_force_src2_zero~q ),
	.datad(\R_ctrl_unsigned_lo_imm16~q ),
	.cin(gnd),
	.combout(\R_src2_hi[15]~2_combout ),
	.cout());
defparam \R_src2_hi[15]~2 .lut_mask = 16'hAFFF;
defparam \R_src2_hi[15]~2 .sum_lutc_input = "datac";

dffeas \E_src2[31] (
	.clk(clk_clk),
	.d(\R_src2_hi[15]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[31]~q ),
	.prn(vcc));
defparam \E_src2[31] .is_wysiwyg = "true";
defparam \E_src2[31] .power_up = "low";

cyclone10lp_lcell_comb \E_invert_arith_src_msb~0 (
	.dataa(\Equal0~9_combout ),
	.datab(\Equal62~0_combout ),
	.datac(\D_iw[14]~q ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\E_invert_arith_src_msb~0_combout ),
	.cout());
defparam \E_invert_arith_src_msb~0 .lut_mask = 16'hEFFE;
defparam \E_invert_arith_src_msb~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_invert_arith_src_msb~1 (
	.dataa(\R_valid~q ),
	.datab(\E_invert_arith_src_msb~0_combout ),
	.datac(\D_iw[5]~q ),
	.datad(\D_ctrl_alu_subtract~2_combout ),
	.cin(gnd),
	.combout(\E_invert_arith_src_msb~1_combout ),
	.cout());
defparam \E_invert_arith_src_msb~1 .lut_mask = 16'hEFFF;
defparam \E_invert_arith_src_msb~1 .sum_lutc_input = "datac";

dffeas E_invert_arith_src_msb(
	.clk(clk_clk),
	.d(\E_invert_arith_src_msb~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_invert_arith_src_msb~q ),
	.prn(vcc));
defparam E_invert_arith_src_msb.is_wysiwyg = "true";
defparam E_invert_arith_src_msb.power_up = "low";

cyclone10lp_lcell_comb \Add1~53 (
	.dataa(\E_alu_sub~q ),
	.datab(\E_src2[31]~q ),
	.datac(\E_invert_arith_src_msb~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add1~53_combout ),
	.cout());
defparam \Add1~53 .lut_mask = 16'h9696;
defparam \Add1~53 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_arith_src1[31] (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_invert_arith_src_msb~q ),
	.datad(\E_src1[31]~q ),
	.cin(gnd),
	.combout(\E_arith_src1[31]~combout ),
	.cout());
defparam \E_arith_src1[31] .lut_mask = 16'h0FF0;
defparam \E_arith_src1[31] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_src2[30]~1 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[30]~1_combout ),
	.cout());
defparam \E_src2[30]~1 .lut_mask = 16'hAACC;
defparam \E_src2[30]~1 .sum_lutc_input = "datac";

dffeas \E_src2[30] (
	.clk(clk_clk),
	.d(\E_src2[30]~1_combout ),
	.asdata(\D_iw[20]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[30]~q ),
	.prn(vcc));
defparam \E_src2[30] .is_wysiwyg = "true";
defparam \E_src2[30] .power_up = "low";

cyclone10lp_lcell_comb \Add1~54 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[30]~q ),
	.cin(gnd),
	.combout(\Add1~54_combout ),
	.cout());
defparam \Add1~54 .lut_mask = 16'h0FF0;
defparam \Add1~54 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_src2[29]~14 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[29]~14_combout ),
	.cout());
defparam \E_src2[29]~14 .lut_mask = 16'hAACC;
defparam \E_src2[29]~14 .sum_lutc_input = "datac";

dffeas \E_src2[29] (
	.clk(clk_clk),
	.d(\E_src2[29]~14_combout ),
	.asdata(\D_iw[19]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[29]~q ),
	.prn(vcc));
defparam \E_src2[29] .is_wysiwyg = "true";
defparam \E_src2[29] .power_up = "low";

cyclone10lp_lcell_comb \Add1~55 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[29]~q ),
	.cin(gnd),
	.combout(\Add1~55_combout ),
	.cout());
defparam \Add1~55 .lut_mask = 16'h0FF0;
defparam \Add1~55 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_src2[28]~2 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[28]~2_combout ),
	.cout());
defparam \E_src2[28]~2 .lut_mask = 16'hAACC;
defparam \E_src2[28]~2 .sum_lutc_input = "datac";

dffeas \E_src2[28] (
	.clk(clk_clk),
	.d(\E_src2[28]~2_combout ),
	.asdata(\D_iw[18]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[28]~q ),
	.prn(vcc));
defparam \E_src2[28] .is_wysiwyg = "true";
defparam \E_src2[28] .power_up = "low";

cyclone10lp_lcell_comb \Add1~56 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[28]~q ),
	.cin(gnd),
	.combout(\Add1~56_combout ),
	.cout());
defparam \Add1~56 .lut_mask = 16'h0FF0;
defparam \Add1~56 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_src2[27]~3 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[27]~3_combout ),
	.cout());
defparam \E_src2[27]~3 .lut_mask = 16'hAACC;
defparam \E_src2[27]~3 .sum_lutc_input = "datac";

dffeas \E_src2[27] (
	.clk(clk_clk),
	.d(\E_src2[27]~3_combout ),
	.asdata(\D_iw[17]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[27]~q ),
	.prn(vcc));
defparam \E_src2[27] .is_wysiwyg = "true";
defparam \E_src2[27] .power_up = "low";

cyclone10lp_lcell_comb \Add1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[27]~q ),
	.cin(gnd),
	.combout(\Add1~57_combout ),
	.cout());
defparam \Add1~57 .lut_mask = 16'h0FF0;
defparam \Add1~57 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_src2[26]~4 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[26]~4_combout ),
	.cout());
defparam \E_src2[26]~4 .lut_mask = 16'hAACC;
defparam \E_src2[26]~4 .sum_lutc_input = "datac";

dffeas \E_src2[26] (
	.clk(clk_clk),
	.d(\E_src2[26]~4_combout ),
	.asdata(\D_iw[16]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[26]~q ),
	.prn(vcc));
defparam \E_src2[26] .is_wysiwyg = "true";
defparam \E_src2[26] .power_up = "low";

cyclone10lp_lcell_comb \Add1~58 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[26]~q ),
	.cin(gnd),
	.combout(\Add1~58_combout ),
	.cout());
defparam \Add1~58 .lut_mask = 16'h0FF0;
defparam \Add1~58 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_src2[25]~5 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[25]~5_combout ),
	.cout());
defparam \E_src2[25]~5 .lut_mask = 16'hAACC;
defparam \E_src2[25]~5 .sum_lutc_input = "datac";

dffeas \E_src2[25] (
	.clk(clk_clk),
	.d(\E_src2[25]~5_combout ),
	.asdata(\D_iw[15]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[25]~q ),
	.prn(vcc));
defparam \E_src2[25] .is_wysiwyg = "true";
defparam \E_src2[25] .power_up = "low";

cyclone10lp_lcell_comb \Add1~59 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[25]~q ),
	.cin(gnd),
	.combout(\Add1~59_combout ),
	.cout());
defparam \Add1~59 .lut_mask = 16'h0FF0;
defparam \Add1~59 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_src2[24]~6 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[24]~6_combout ),
	.cout());
defparam \E_src2[24]~6 .lut_mask = 16'hAACC;
defparam \E_src2[24]~6 .sum_lutc_input = "datac";

dffeas \E_src2[24] (
	.clk(clk_clk),
	.d(\E_src2[24]~6_combout ),
	.asdata(\D_iw[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[24]~q ),
	.prn(vcc));
defparam \E_src2[24] .is_wysiwyg = "true";
defparam \E_src2[24] .power_up = "low";

cyclone10lp_lcell_comb \Add1~60 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[24]~q ),
	.cin(gnd),
	.combout(\Add1~60_combout ),
	.cout());
defparam \Add1~60 .lut_mask = 16'h0FF0;
defparam \Add1~60 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_src2[23]~7 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[23]~7_combout ),
	.cout());
defparam \E_src2[23]~7 .lut_mask = 16'hAACC;
defparam \E_src2[23]~7 .sum_lutc_input = "datac";

dffeas \E_src2[23] (
	.clk(clk_clk),
	.d(\E_src2[23]~7_combout ),
	.asdata(\D_iw[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[23]~q ),
	.prn(vcc));
defparam \E_src2[23] .is_wysiwyg = "true";
defparam \E_src2[23] .power_up = "low";

cyclone10lp_lcell_comb \Add1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[23]~q ),
	.cin(gnd),
	.combout(\Add1~61_combout ),
	.cout());
defparam \Add1~61 .lut_mask = 16'h0FF0;
defparam \Add1~61 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_src2[22]~8 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[22]~8_combout ),
	.cout());
defparam \E_src2[22]~8 .lut_mask = 16'hAACC;
defparam \E_src2[22]~8 .sum_lutc_input = "datac";

dffeas \E_src2[22] (
	.clk(clk_clk),
	.d(\E_src2[22]~8_combout ),
	.asdata(\D_iw[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[22]~q ),
	.prn(vcc));
defparam \E_src2[22] .is_wysiwyg = "true";
defparam \E_src2[22] .power_up = "low";

cyclone10lp_lcell_comb \Add1~62 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[22]~q ),
	.cin(gnd),
	.combout(\Add1~62_combout ),
	.cout());
defparam \Add1~62 .lut_mask = 16'h0FF0;
defparam \Add1~62 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_src2[21]~9 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[21]~9_combout ),
	.cout());
defparam \E_src2[21]~9 .lut_mask = 16'hAACC;
defparam \E_src2[21]~9 .sum_lutc_input = "datac";

dffeas \E_src2[21] (
	.clk(clk_clk),
	.d(\E_src2[21]~9_combout ),
	.asdata(\D_iw[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[21]~q ),
	.prn(vcc));
defparam \E_src2[21] .is_wysiwyg = "true";
defparam \E_src2[21] .power_up = "low";

cyclone10lp_lcell_comb \Add1~63 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[21]~q ),
	.cin(gnd),
	.combout(\Add1~63_combout ),
	.cout());
defparam \Add1~63 .lut_mask = 16'h0FF0;
defparam \Add1~63 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_src2[20]~10 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[20]~10_combout ),
	.cout());
defparam \E_src2[20]~10 .lut_mask = 16'hAACC;
defparam \E_src2[20]~10 .sum_lutc_input = "datac";

dffeas \E_src2[20] (
	.clk(clk_clk),
	.d(\E_src2[20]~10_combout ),
	.asdata(\D_iw[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[20]~q ),
	.prn(vcc));
defparam \E_src2[20] .is_wysiwyg = "true";
defparam \E_src2[20] .power_up = "low";

cyclone10lp_lcell_comb \Add1~64 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[20]~q ),
	.cin(gnd),
	.combout(\Add1~64_combout ),
	.cout());
defparam \Add1~64 .lut_mask = 16'h0FF0;
defparam \Add1~64 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_src2[19]~11 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[19]~11_combout ),
	.cout());
defparam \E_src2[19]~11 .lut_mask = 16'hAACC;
defparam \E_src2[19]~11 .sum_lutc_input = "datac";

dffeas \E_src2[19] (
	.clk(clk_clk),
	.d(\E_src2[19]~11_combout ),
	.asdata(\D_iw[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[19]~q ),
	.prn(vcc));
defparam \E_src2[19] .is_wysiwyg = "true";
defparam \E_src2[19] .power_up = "low";

cyclone10lp_lcell_comb \Add1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[19]~q ),
	.cin(gnd),
	.combout(\Add1~65_combout ),
	.cout());
defparam \Add1~65 .lut_mask = 16'h0FF0;
defparam \Add1~65 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_src2[18]~12 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[18]~12_combout ),
	.cout());
defparam \E_src2[18]~12 .lut_mask = 16'hAACC;
defparam \E_src2[18]~12 .sum_lutc_input = "datac";

dffeas \E_src2[18] (
	.clk(clk_clk),
	.d(\E_src2[18]~12_combout ),
	.asdata(\D_iw[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[18]~q ),
	.prn(vcc));
defparam \E_src2[18] .is_wysiwyg = "true";
defparam \E_src2[18] .power_up = "low";

cyclone10lp_lcell_comb \Add1~66 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[18]~q ),
	.cin(gnd),
	.combout(\Add1~66_combout ),
	.cout());
defparam \Add1~66 .lut_mask = 16'h0FF0;
defparam \Add1~66 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_src2[17]~13 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[17]~13_combout ),
	.cout());
defparam \E_src2[17]~13 .lut_mask = 16'hAACC;
defparam \E_src2[17]~13 .sum_lutc_input = "datac";

dffeas \E_src2[17] (
	.clk(clk_clk),
	.d(\E_src2[17]~13_combout ),
	.asdata(\D_iw[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[17]~q ),
	.prn(vcc));
defparam \E_src2[17] .is_wysiwyg = "true";
defparam \E_src2[17] .power_up = "low";

cyclone10lp_lcell_comb \Add1~67 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[17]~q ),
	.cin(gnd),
	.combout(\Add1~67_combout ),
	.cout());
defparam \Add1~67 .lut_mask = 16'h0FF0;
defparam \Add1~67 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Add1~98 (
	.dataa(\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add1~97 ),
	.combout(\Add1~98_combout ),
	.cout());
defparam \Add1~98 .lut_mask = 16'h5A5A;
defparam \Add1~98 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Equal127~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_logic_result[16]~1_combout ),
	.datad(\E_logic_result[15]~2_combout ),
	.cin(gnd),
	.combout(\Equal127~0_combout ),
	.cout());
defparam \Equal127~0 .lut_mask = 16'h0FFF;
defparam \Equal127~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal127~1 (
	.dataa(\E_logic_result[12]~5_combout ),
	.datab(\E_logic_result[11]~6_combout ),
	.datac(\E_logic_result[10]~7_combout ),
	.datad(\E_logic_result[9]~8_combout ),
	.cin(gnd),
	.combout(\Equal127~1_combout ),
	.cout());
defparam \Equal127~1 .lut_mask = 16'h7FFF;
defparam \Equal127~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal127~2 (
	.dataa(\Equal127~0_combout ),
	.datab(\Equal127~1_combout ),
	.datac(\E_logic_result[14]~3_combout ),
	.datad(\E_logic_result[13]~4_combout ),
	.cin(gnd),
	.combout(\Equal127~2_combout ),
	.cout());
defparam \Equal127~2 .lut_mask = 16'hEFFF;
defparam \Equal127~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal127~3 (
	.dataa(\E_logic_result[5]~11_combout ),
	.datab(\E_logic_result[6]~12_combout ),
	.datac(\E_logic_result[7]~0_combout ),
	.datad(\E_logic_result[8]~9_combout ),
	.cin(gnd),
	.combout(\Equal127~3_combout ),
	.cout());
defparam \Equal127~3 .lut_mask = 16'h7FFF;
defparam \Equal127~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_logic_result[31]~15 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[31]~q ),
	.datac(\E_src1[31]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[31]~15_combout ),
	.cout());
defparam \E_logic_result[31]~15 .lut_mask = 16'h6996;
defparam \E_logic_result[31]~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal127~4 (
	.dataa(\E_logic_result[4]~10_combout ),
	.datab(\E_logic_result[2]~13_combout ),
	.datac(\E_logic_result[3]~14_combout ),
	.datad(\E_logic_result[31]~15_combout ),
	.cin(gnd),
	.combout(\Equal127~4_combout ),
	.cout());
defparam \Equal127~4 .lut_mask = 16'h7FFF;
defparam \Equal127~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_logic_result[30]~16 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[30]~q ),
	.datac(\E_src1[30]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[30]~16_combout ),
	.cout());
defparam \E_logic_result[30]~16 .lut_mask = 16'h6996;
defparam \E_logic_result[30]~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_logic_result[28]~17 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[28]~q ),
	.datac(\E_src1[28]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[28]~17_combout ),
	.cout());
defparam \E_logic_result[28]~17 .lut_mask = 16'h6996;
defparam \E_logic_result[28]~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_logic_result[27]~18 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[27]~q ),
	.datac(\E_src1[27]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[27]~18_combout ),
	.cout());
defparam \E_logic_result[27]~18 .lut_mask = 16'h6996;
defparam \E_logic_result[27]~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_logic_result[26]~19 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[26]~q ),
	.datac(\E_src1[26]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[26]~19_combout ),
	.cout());
defparam \E_logic_result[26]~19 .lut_mask = 16'h6996;
defparam \E_logic_result[26]~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal127~5 (
	.dataa(\E_logic_result[30]~16_combout ),
	.datab(\E_logic_result[28]~17_combout ),
	.datac(\E_logic_result[27]~18_combout ),
	.datad(\E_logic_result[26]~19_combout ),
	.cin(gnd),
	.combout(\Equal127~5_combout ),
	.cout());
defparam \Equal127~5 .lut_mask = 16'h7FFF;
defparam \Equal127~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_logic_result[25]~20 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[25]~q ),
	.datac(\E_src1[25]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[25]~20_combout ),
	.cout());
defparam \E_logic_result[25]~20 .lut_mask = 16'h6996;
defparam \E_logic_result[25]~20 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_logic_result[24]~21 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[24]~q ),
	.datac(\E_src1[24]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[24]~21_combout ),
	.cout());
defparam \E_logic_result[24]~21 .lut_mask = 16'h6996;
defparam \E_logic_result[24]~21 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_logic_result[23]~22 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[23]~q ),
	.datac(\E_src1[23]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[23]~22_combout ),
	.cout());
defparam \E_logic_result[23]~22 .lut_mask = 16'h6996;
defparam \E_logic_result[23]~22 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_logic_result[22]~23 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[22]~q ),
	.datac(\E_src1[22]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[22]~23_combout ),
	.cout());
defparam \E_logic_result[22]~23 .lut_mask = 16'h6996;
defparam \E_logic_result[22]~23 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal127~6 (
	.dataa(\E_logic_result[25]~20_combout ),
	.datab(\E_logic_result[24]~21_combout ),
	.datac(\E_logic_result[23]~22_combout ),
	.datad(\E_logic_result[22]~23_combout ),
	.cin(gnd),
	.combout(\Equal127~6_combout ),
	.cout());
defparam \Equal127~6 .lut_mask = 16'h7FFF;
defparam \Equal127~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_logic_result[21]~24 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[21]~q ),
	.datac(\E_src1[21]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[21]~24_combout ),
	.cout());
defparam \E_logic_result[21]~24 .lut_mask = 16'h6996;
defparam \E_logic_result[21]~24 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_logic_result[20]~25 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[20]~q ),
	.datac(\E_src1[20]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[20]~25_combout ),
	.cout());
defparam \E_logic_result[20]~25 .lut_mask = 16'h6996;
defparam \E_logic_result[20]~25 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_logic_result[19]~26 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[19]~q ),
	.datac(\E_src1[19]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[19]~26_combout ),
	.cout());
defparam \E_logic_result[19]~26 .lut_mask = 16'h6996;
defparam \E_logic_result[19]~26 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_logic_result[18]~27 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[18]~q ),
	.datac(\E_src1[18]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[18]~27_combout ),
	.cout());
defparam \E_logic_result[18]~27 .lut_mask = 16'h6996;
defparam \E_logic_result[18]~27 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal127~7 (
	.dataa(\E_logic_result[21]~24_combout ),
	.datab(\E_logic_result[20]~25_combout ),
	.datac(\E_logic_result[19]~26_combout ),
	.datad(\E_logic_result[18]~27_combout ),
	.cin(gnd),
	.combout(\Equal127~7_combout ),
	.cout());
defparam \Equal127~7 .lut_mask = 16'h7FFF;
defparam \Equal127~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_logic_result[17]~28 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[17]~q ),
	.datac(\E_src1[17]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[17]~28_combout ),
	.cout());
defparam \E_logic_result[17]~28 .lut_mask = 16'h6996;
defparam \E_logic_result[17]~28 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_logic_result[1]~29 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[1]~q ),
	.datac(\E_src1[1]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[1]~29_combout ),
	.cout());
defparam \E_logic_result[1]~29 .lut_mask = 16'h6996;
defparam \E_logic_result[1]~29 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_logic_result[0]~30 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[0]~q ),
	.datac(\E_src1[0]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[0]~30_combout ),
	.cout());
defparam \E_logic_result[0]~30 .lut_mask = 16'h6996;
defparam \E_logic_result[0]~30 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_logic_result[29]~31 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[29]~q ),
	.datac(\E_src1[29]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[29]~31_combout ),
	.cout());
defparam \E_logic_result[29]~31 .lut_mask = 16'h6996;
defparam \E_logic_result[29]~31 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal127~8 (
	.dataa(\E_logic_result[17]~28_combout ),
	.datab(\E_logic_result[1]~29_combout ),
	.datac(\E_logic_result[0]~30_combout ),
	.datad(\E_logic_result[29]~31_combout ),
	.cin(gnd),
	.combout(\Equal127~8_combout ),
	.cout());
defparam \Equal127~8 .lut_mask = 16'h7FFF;
defparam \Equal127~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal127~9 (
	.dataa(\Equal127~5_combout ),
	.datab(\Equal127~6_combout ),
	.datac(\Equal127~7_combout ),
	.datad(\Equal127~8_combout ),
	.cin(gnd),
	.combout(\Equal127~9_combout ),
	.cout());
defparam \Equal127~9 .lut_mask = 16'hFFFE;
defparam \Equal127~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal127~10 (
	.dataa(\Equal127~2_combout ),
	.datab(\Equal127~3_combout ),
	.datac(\Equal127~4_combout ),
	.datad(\Equal127~9_combout ),
	.cin(gnd),
	.combout(\Equal127~10_combout ),
	.cout());
defparam \Equal127~10 .lut_mask = 16'hFFFE;
defparam \Equal127~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \D_logic_op_raw[0]~1 (
	.dataa(\D_iw[14]~q ),
	.datab(\D_iw[3]~q ),
	.datac(\Equal0~4_combout ),
	.datad(\Equal0~5_combout ),
	.cin(gnd),
	.combout(\D_logic_op_raw[0]~1_combout ),
	.cout());
defparam \D_logic_op_raw[0]~1 .lut_mask = 16'hEFFE;
defparam \D_logic_op_raw[0]~1 .sum_lutc_input = "datac";

dffeas \R_compare_op[0] (
	.clk(clk_clk),
	.d(\D_logic_op_raw[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_compare_op[0]~q ),
	.prn(vcc));
defparam \R_compare_op[0] .is_wysiwyg = "true";
defparam \R_compare_op[0] .power_up = "low";

cyclone10lp_lcell_comb \E_cmp_result~0 (
	.dataa(\R_compare_op[1]~q ),
	.datab(\Add1~98_combout ),
	.datac(\Equal127~10_combout ),
	.datad(\R_compare_op[0]~q ),
	.cin(gnd),
	.combout(\E_cmp_result~0_combout ),
	.cout());
defparam \E_cmp_result~0 .lut_mask = 16'h6996;
defparam \E_cmp_result~0 .sum_lutc_input = "datac";

dffeas W_cmp_result(
	.clk(clk_clk),
	.d(\E_cmp_result~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_cmp_result~q ),
	.prn(vcc));
defparam W_cmp_result.is_wysiwyg = "true";
defparam W_cmp_result.power_up = "low";

cyclone10lp_lcell_comb \F_pc_sel_nxt~0 (
	.dataa(\R_ctrl_uncond_cti_non_br~q ),
	.datab(\R_ctrl_br_uncond~q ),
	.datac(\W_cmp_result~q ),
	.datad(\R_ctrl_br~q ),
	.cin(gnd),
	.combout(\F_pc_sel_nxt~0_combout ),
	.cout());
defparam \F_pc_sel_nxt~0 .lut_mask = 16'hFFFE;
defparam \F_pc_sel_nxt~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_pc_sel_nxt.10~0 (
	.dataa(\F_pc_sel_nxt~0_combout ),
	.datab(gnd),
	.datac(\R_ctrl_exception~q ),
	.datad(\R_ctrl_break~q ),
	.cin(gnd),
	.combout(\F_pc_sel_nxt.10~0_combout ),
	.cout());
defparam \F_pc_sel_nxt.10~0 .lut_mask = 16'hAFFF;
defparam \F_pc_sel_nxt.10~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_pc_no_crst_nxt[5]~0 (
	.dataa(\Add1~24_combout ),
	.datab(\F_pc_plus_one[5]~10_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[5]~0_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[5]~0 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[5]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_pc_no_crst_nxt[14]~1 (
	.dataa(\R_ctrl_break~q ),
	.datab(\F_pc_plus_one[14]~28_combout ),
	.datac(gnd),
	.datad(\F_pc_sel_nxt~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[14]~1_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[14]~1 .lut_mask = 16'hEEFF;
defparam \F_pc_no_crst_nxt[14]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_pc_no_crst_nxt[14]~2 (
	.dataa(\F_pc_no_crst_nxt[14]~1_combout ),
	.datab(\F_pc_sel_nxt~0_combout ),
	.datac(\Add1~51_combout ),
	.datad(\R_ctrl_exception~q ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[14]~2_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[14]~2 .lut_mask = 16'hFEFF;
defparam \F_pc_no_crst_nxt[14]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_pc_no_crst_nxt[13]~3 (
	.dataa(\F_pc_plus_one[13]~26_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\R_ctrl_break~q ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[13]~3_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[13]~3 .lut_mask = 16'hAAFF;
defparam \F_pc_no_crst_nxt[13]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_pc_no_crst_nxt[13]~4 (
	.dataa(\R_ctrl_exception~q ),
	.datab(\Add1~49_combout ),
	.datac(\F_pc_no_crst_nxt[13]~3_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[13]~4_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[13]~4 .lut_mask = 16'h5F3F;
defparam \F_pc_no_crst_nxt[13]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_pc_no_crst_nxt[12]~5 (
	.dataa(\Add1~47_combout ),
	.datab(\F_pc_plus_one[12]~24_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[12]~5_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[12]~5 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[12]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_pc_no_crst_nxt[11]~6 (
	.dataa(\Add1~45_combout ),
	.datab(\F_pc_plus_one[11]~22_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[11]~6_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[11]~6 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[11]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_pc_no_crst_nxt[10]~7 (
	.dataa(\Add1~43_combout ),
	.datab(\F_pc_plus_one[10]~20_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[10]~7_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[10]~7 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[10]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_pc_no_crst_nxt[9]~8 (
	.dataa(\F_pc_plus_one[9]~18_combout ),
	.datab(\Add1~41_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[9]~8_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[9]~8 .lut_mask = 16'hEFFE;
defparam \F_pc_no_crst_nxt[9]~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_pc_no_crst_nxt[9]~9 (
	.dataa(\R_ctrl_break~q ),
	.datab(\F_pc_no_crst_nxt[9]~8_combout ),
	.datac(gnd),
	.datad(\R_ctrl_exception~q ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[9]~9_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[9]~9 .lut_mask = 16'hEEFF;
defparam \F_pc_no_crst_nxt[9]~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_pc_no_crst_nxt[8]~10 (
	.dataa(\Add1~39_combout ),
	.datab(\F_pc_plus_one[8]~16_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[8]~10_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[8]~10 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[8]~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_pc_no_crst_nxt[7]~11 (
	.dataa(\Add1~37_combout ),
	.datab(\F_pc_plus_one[7]~14_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[7]~11_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[7]~11 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[7]~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_pc_no_crst_nxt[6]~12 (
	.dataa(\Add1~35_combout ),
	.datab(\F_pc_plus_one[6]~12_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[6]~12_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[6]~12 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[6]~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_pc_no_crst_nxt[2]~13 (
	.dataa(\Add1~18_combout ),
	.datab(\F_pc_plus_one[2]~4_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[2]~13_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[2]~13 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[2]~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_pc_no_crst_nxt[3]~14 (
	.dataa(\F_pc_sel_nxt.10~1_combout ),
	.datab(\Add1~20_combout ),
	.datac(\F_pc_plus_one[3]~6_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[3]~14_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[3]~14 .lut_mask = 16'hFAFC;
defparam \F_pc_no_crst_nxt[3]~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_pc_no_crst_nxt[4]~15 (
	.dataa(\Add1~22_combout ),
	.datab(\F_pc_plus_one[4]~8_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[4]~15_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[4]~15 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[4]~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb d_read_nxt(
	.dataa(d_read1),
	.datab(\E_new_inst~q ),
	.datac(\R_ctrl_ld~q ),
	.datad(WideOr12),
	.cin(gnd),
	.combout(\d_read_nxt~combout ),
	.cout());
defparam d_read_nxt.lut_mask = 16'hFFFE;
defparam d_read_nxt.sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_pc_no_crst_nxt[1]~16 (
	.dataa(\Add1~16_combout ),
	.datab(\F_pc_plus_one[1]~2_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[1]~16_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[1]~16 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[1]~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \F_pc_no_crst_nxt[0]~17 (
	.dataa(\Add1~14_combout ),
	.datab(\F_pc_plus_one[0]~0_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[0]~17_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[0]~17 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[0]~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_st_data[9]~0 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[9]~0_combout ),
	.cout());
defparam \E_st_data[9]~0 .lut_mask = 16'hEFFE;
defparam \E_st_data[9]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \hbreak_enabled~0 (
	.dataa(\D_op_cmpge~0_combout ),
	.datab(\Equal62~4_combout ),
	.datac(hbreak_enabled1),
	.datad(\R_ctrl_break~q ),
	.cin(gnd),
	.combout(\hbreak_enabled~0_combout ),
	.cout());
defparam \hbreak_enabled~0 .lut_mask = 16'hFFF7;
defparam \hbreak_enabled~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_mem_byte_en[0]~0 (
	.dataa(\D_ctrl_mem16~1_combout ),
	.datab(\D_ctrl_mem8~1_combout ),
	.datac(\Add1~10_combout ),
	.datad(\Add1~12_combout ),
	.cin(gnd),
	.combout(\E_mem_byte_en[0]~0_combout ),
	.cout());
defparam \E_mem_byte_en[0]~0 .lut_mask = 16'h6FFF;
defparam \E_mem_byte_en[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \d_byteenable[2]~0 (
	.dataa(\D_ctrl_mem16~0_combout ),
	.datab(\D_ctrl_mem8~0_combout ),
	.datac(gnd),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\d_byteenable[2]~0_combout ),
	.cout());
defparam \d_byteenable[2]~0 .lut_mask = 16'hEEFF;
defparam \d_byteenable[2]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_st_data[22]~1 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.datac(gnd),
	.datad(\d_byteenable[2]~0_combout ),
	.cin(gnd),
	.combout(\E_st_data[22]~1_combout ),
	.cout());
defparam \E_st_data[22]~1 .lut_mask = 16'hAACC;
defparam \E_st_data[22]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_mem_byte_en[2]~1 (
	.dataa(\D_ctrl_mem16~1_combout ),
	.datab(\Add1~12_combout ),
	.datac(\D_ctrl_mem8~1_combout ),
	.datad(\Add1~10_combout ),
	.cin(gnd),
	.combout(\E_mem_byte_en[2]~1_combout ),
	.cout());
defparam \E_mem_byte_en[2]~1 .lut_mask = 16'hDEFF;
defparam \E_mem_byte_en[2]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_st_data[23]~2 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.datac(gnd),
	.datad(\d_byteenable[2]~0_combout ),
	.cin(gnd),
	.combout(\E_st_data[23]~2_combout ),
	.cout());
defparam \E_st_data[23]~2 .lut_mask = 16'hAACC;
defparam \E_st_data[23]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_mem_byte_en[3]~2 (
	.dataa(\D_ctrl_mem16~1_combout ),
	.datab(\Add1~12_combout ),
	.datac(\Add1~10_combout ),
	.datad(\D_ctrl_mem8~1_combout ),
	.cin(gnd),
	.combout(\E_mem_byte_en[3]~2_combout ),
	.cout());
defparam \E_mem_byte_en[3]~2 .lut_mask = 16'hFDFE;
defparam \E_mem_byte_en[3]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_st_data[14]~3 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[14]~3_combout ),
	.cout());
defparam \E_st_data[14]~3 .lut_mask = 16'hEFFE;
defparam \E_st_data[14]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_mem_byte_en[1]~3 (
	.dataa(\D_ctrl_mem16~1_combout ),
	.datab(\D_ctrl_mem8~1_combout ),
	.datac(\Add1~10_combout ),
	.datad(\Add1~12_combout ),
	.cin(gnd),
	.combout(\E_mem_byte_en[1]~3_combout ),
	.cout());
defparam \E_mem_byte_en[1]~3 .lut_mask = 16'hF6FF;
defparam \E_mem_byte_en[1]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_st_data[15]~4 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[15]~4_combout ),
	.cout());
defparam \E_st_data[15]~4 .lut_mask = 16'hEFFE;
defparam \E_st_data[15]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_st_data[11]~5 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[11]~5_combout ),
	.cout());
defparam \E_st_data[11]~5 .lut_mask = 16'hEFFE;
defparam \E_st_data[11]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_st_data[13]~6 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[13]~6_combout ),
	.cout());
defparam \E_st_data[13]~6 .lut_mask = 16'hEFFE;
defparam \E_st_data[13]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_st_data[16]~7 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.datac(gnd),
	.datad(\d_byteenable[2]~0_combout ),
	.cin(gnd),
	.combout(\E_st_data[16]~7_combout ),
	.cout());
defparam \E_st_data[16]~7 .lut_mask = 16'hAACC;
defparam \E_st_data[16]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_st_data[12]~8 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[12]~8_combout ),
	.cout());
defparam \E_st_data[12]~8 .lut_mask = 16'hEFFE;
defparam \E_st_data[12]~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_st_data[10]~9 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[10]~9_combout ),
	.cout());
defparam \E_st_data[10]~9 .lut_mask = 16'hEFFE;
defparam \E_st_data[10]~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_st_data[8]~10 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[8]~10_combout ),
	.cout());
defparam \E_st_data[8]~10 .lut_mask = 16'hEFFE;
defparam \E_st_data[8]~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_st_data[21]~11 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.datac(gnd),
	.datad(\d_byteenable[2]~0_combout ),
	.cin(gnd),
	.combout(\E_st_data[21]~11_combout ),
	.cout());
defparam \E_st_data[21]~11 .lut_mask = 16'hAACC;
defparam \E_st_data[21]~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_st_data[20]~12 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ),
	.datac(gnd),
	.datad(\d_byteenable[2]~0_combout ),
	.cin(gnd),
	.combout(\E_st_data[20]~12_combout ),
	.cout());
defparam \E_st_data[20]~12 .lut_mask = 16'hAACC;
defparam \E_st_data[20]~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_st_data[19]~13 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ),
	.datac(gnd),
	.datad(\d_byteenable[2]~0_combout ),
	.cin(gnd),
	.combout(\E_st_data[19]~13_combout ),
	.cout());
defparam \E_st_data[19]~13 .lut_mask = 16'hAACC;
defparam \E_st_data[19]~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_st_data[18]~14 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.datac(gnd),
	.datad(\d_byteenable[2]~0_combout ),
	.cin(gnd),
	.combout(\E_st_data[18]~14_combout ),
	.cout());
defparam \E_st_data[18]~14 .lut_mask = 16'hAACC;
defparam \E_st_data[18]~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \E_st_data[17]~15 (
	.dataa(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.datab(\processor_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.datac(gnd),
	.datad(\d_byteenable[2]~0_combout ),
	.cin(gnd),
	.combout(\E_st_data[17]~15_combout ),
	.cout());
defparam \E_st_data[17]~15 .lut_mask = 16'hAACC;
defparam \E_st_data[17]~15 .sum_lutc_input = "datac";

endmodule

module processor_processor_nios2_gen2_0_cpu_nios2_oci (
	sr_0,
	jtag_break,
	readdata_0,
	readdata_1,
	readdata_3,
	readdata_2,
	ir_out_0,
	ir_out_1,
	r_sync_rst,
	saved_grant_0,
	waitrequest,
	mem_used_1,
	uav_write,
	WideOr1,
	rf_source_valid,
	hbreak_enabled,
	address_nxt,
	r_early_rst,
	oci_ienable_0,
	oci_ienable_1,
	oci_single_step_mode,
	readdata_22,
	readdata_23,
	readdata_24,
	readdata_25,
	readdata_26,
	readdata_4,
	readdata_5,
	readdata_14,
	readdata_15,
	readdata_11,
	readdata_13,
	readdata_16,
	readdata_12,
	readdata_10,
	readdata_9,
	readdata_8,
	readdata_7,
	readdata_6,
	readdata_21,
	readdata_20,
	readdata_19,
	readdata_18,
	readdata_17,
	debugaccess_nxt,
	writedata_nxt,
	byteenable_nxt,
	readdata_27,
	readdata_28,
	readdata_29,
	readdata_30,
	readdata_31,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	sr_0;
output 	jtag_break;
output 	readdata_0;
output 	readdata_1;
output 	readdata_3;
output 	readdata_2;
output 	ir_out_0;
output 	ir_out_1;
input 	r_sync_rst;
input 	saved_grant_0;
output 	waitrequest;
input 	mem_used_1;
input 	uav_write;
input 	WideOr1;
input 	rf_source_valid;
input 	hbreak_enabled;
input 	[8:0] address_nxt;
input 	r_early_rst;
output 	oci_ienable_0;
output 	oci_ienable_1;
output 	oci_single_step_mode;
output 	readdata_22;
output 	readdata_23;
output 	readdata_24;
output 	readdata_25;
output 	readdata_26;
output 	readdata_4;
output 	readdata_5;
output 	readdata_14;
output 	readdata_15;
output 	readdata_11;
output 	readdata_13;
output 	readdata_16;
output 	readdata_12;
output 	readdata_10;
output 	readdata_9;
output 	readdata_8;
output 	readdata_7;
output 	readdata_6;
output 	readdata_21;
output 	readdata_20;
output 	readdata_19;
output 	readdata_18;
output 	readdata_17;
input 	debugaccess_nxt;
input 	[31:0] writedata_nxt;
input 	[3:0] byteenable_nxt;
output 	readdata_27;
output 	readdata_28;
output 	readdata_29;
output 	readdata_30;
output 	readdata_31;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[0]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[4]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[29]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[5]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[15]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[12]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[8]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[18]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[0]~q ;
wire \write~q ;
wire \read~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[1]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[1]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[0]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[36]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[37]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|ir[0]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|ir[1]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|enable_action_strobe~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[3]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[35]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|take_action_ocimem_b~combout ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|take_action_ocimem_a~0_combout ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_debug|monitor_ready~q ;
wire \write~0_combout ;
wire \write~1_combout ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[17]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|take_action_ocimem_a~1_combout ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[34]~q ;
wire \read~0_combout ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[2]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[2]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[1]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[4]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[26]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[28]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[27]~q ;
wire \debugaccess~q ;
wire \writedata[0]~q ;
wire \address[0]~q ;
wire \address[1]~q ;
wire \address[2]~q ;
wire \address[3]~q ;
wire \address[4]~q ;
wire \address[5]~q ;
wire \address[6]~q ;
wire \address[7]~q ;
wire \byteenable[0]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal0~2_combout ;
wire \the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|take_action_ocireg~0_combout ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[25]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[21]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[20]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|take_action_ocimem_a~combout ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[33]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[32]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[31]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[30]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[29]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[3]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[3]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[2]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[5]~q ;
wire \writedata[1]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_debug|monitor_error~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[19]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[18]~q ;
wire \writedata[3]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_debug|monitor_go~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[16]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[16]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[4]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[6]~q ;
wire \writedata[2]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[25]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[25]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[27]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[27]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[26]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[26]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[24]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[24]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[20]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[20]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[19]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[19]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[22]~q ;
wire \writedata[22]~q ;
wire \byteenable[2]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[23]~q ;
wire \writedata[23]~q ;
wire \writedata[24]~q ;
wire \byteenable[3]~q ;
wire \writedata[25]~q ;
wire \writedata[26]~q ;
wire \writedata[4]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[23]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[17]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[17]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[16]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_debug|resetlatch~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[31]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[31]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[30]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[30]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[29]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[28]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[28]~q ;
wire \writedata[5]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[14]~q ;
wire \writedata[14]~q ;
wire \byteenable[1]~q ;
wire \writedata[15]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[11]~q ;
wire \writedata[11]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[13]~q ;
wire \writedata[13]~q ;
wire \writedata[16]~q ;
wire \writedata[12]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[10]~q ;
wire \writedata[10]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[9]~q ;
wire \writedata[9]~q ;
wire \writedata[8]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[7]~q ;
wire \writedata[7]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[6]~q ;
wire \writedata[6]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[21]~q ;
wire \writedata[21]~q ;
wire \writedata[20]~q ;
wire \writedata[19]~q ;
wire \writedata[18]~q ;
wire \writedata[17]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[5]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[7]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[24]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[18]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[21]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[22]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[8]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[14]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[15]~q ;
wire \writedata[27]~q ;
wire \writedata[28]~q ;
wire \writedata[29]~q ;
wire \writedata[30]~q ;
wire \writedata[31]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[13]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[12]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[11]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[10]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[9]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[6]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[22]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[15]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[7]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[23]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[13]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[14]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[12]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[11]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[10]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[9]~q ;
wire \the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[8]~q ;
wire \readdata~0_combout ;
wire \address[8]~q ;
wire \readdata~6_combout ;
wire \readdata~8_combout ;
wire \readdata~9_combout ;
wire \readdata~1_combout ;
wire \readdata~2_combout ;
wire \readdata~3_combout ;
wire \readdata~4_combout ;
wire \readdata~5_combout ;
wire \readdata~7_combout ;
wire \readdata~10_combout ;
wire \readdata~11_combout ;
wire \readdata~12_combout ;
wire \readdata~13_combout ;
wire \readdata~14_combout ;
wire \readdata~15_combout ;
wire \readdata~16_combout ;
wire \readdata~17_combout ;
wire \readdata~18_combout ;
wire \readdata~19_combout ;
wire \readdata~20_combout ;
wire \readdata~21_combout ;
wire \readdata~22_combout ;
wire \readdata~23_combout ;
wire \readdata~24_combout ;
wire \readdata~25_combout ;
wire \readdata~26_combout ;
wire \readdata~27_combout ;
wire \readdata~28_combout ;
wire \readdata~29_combout ;
wire \readdata~30_combout ;
wire \readdata~31_combout ;


processor_processor_nios2_gen2_0_cpu_nios2_oci_break the_processor_nios2_gen2_0_cpu_nios2_oci_break(
	.break_readreg_0(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[0]~q ),
	.break_readreg_1(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[1]~q ),
	.jdo_0(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[0]~q ),
	.jdo_36(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[36]~q ),
	.jdo_37(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[37]~q ),
	.ir_0(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|ir[0]~q ),
	.ir_1(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|ir[1]~q ),
	.enable_action_strobe(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|enable_action_strobe~q ),
	.jdo_3(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[3]~q ),
	.jdo_17(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[17]~q ),
	.break_readreg_2(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[2]~q ),
	.jdo_1(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[1]~q ),
	.jdo_4(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[4]~q ),
	.jdo_26(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[26]~q ),
	.jdo_28(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[28]~q ),
	.jdo_27(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[27]~q ),
	.jdo_25(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[25]~q ),
	.jdo_21(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[20]~q ),
	.jdo_31(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[31]~q ),
	.jdo_30(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[30]~q ),
	.jdo_29(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[29]~q ),
	.break_readreg_3(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[3]~q ),
	.jdo_2(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[2]~q ),
	.jdo_5(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[5]~q ),
	.jdo_19(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[18]~q ),
	.break_readreg_16(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[16]~q ),
	.break_readreg_4(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[4]~q ),
	.jdo_6(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[6]~q ),
	.break_readreg_25(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[25]~q ),
	.break_readreg_27(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[27]~q ),
	.break_readreg_26(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[26]~q ),
	.break_readreg_24(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[24]~q ),
	.break_readreg_20(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[20]~q ),
	.break_readreg_19(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[19]~q ),
	.jdo_23(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[23]~q ),
	.break_readreg_17(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[17]~q ),
	.jdo_16(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[16]~q ),
	.break_readreg_31(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[31]~q ),
	.break_readreg_30(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[30]~q ),
	.break_readreg_29(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[29]~q ),
	.break_readreg_28(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[28]~q ),
	.break_readreg_5(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[5]~q ),
	.jdo_7(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[7]~q ),
	.jdo_24(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[24]~q ),
	.break_readreg_18(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[18]~q ),
	.break_readreg_21(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[21]~q ),
	.jdo_22(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[22]~q ),
	.jdo_8(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[8]~q ),
	.jdo_14(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[14]~q ),
	.jdo_15(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[15]~q ),
	.jdo_13(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[13]~q ),
	.jdo_12(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[12]~q ),
	.jdo_11(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[11]~q ),
	.jdo_10(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[10]~q ),
	.jdo_9(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[9]~q ),
	.break_readreg_6(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[6]~q ),
	.break_readreg_22(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[22]~q ),
	.break_readreg_15(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[15]~q ),
	.break_readreg_7(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[7]~q ),
	.break_readreg_23(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[23]~q ),
	.break_readreg_13(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[13]~q ),
	.break_readreg_14(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[14]~q ),
	.break_readreg_12(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[12]~q ),
	.break_readreg_11(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[11]~q ),
	.break_readreg_10(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[10]~q ),
	.break_readreg_9(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[9]~q ),
	.break_readreg_8(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[8]~q ),
	.clk_clk(clk_clk));

processor_processor_nios2_gen2_0_cpu_nios2_oci_debug the_processor_nios2_gen2_0_cpu_nios2_oci_debug(
	.jtag_break1(jtag_break),
	.r_sync_rst(r_sync_rst),
	.monitor_ready1(\the_processor_nios2_gen2_0_cpu_nios2_oci_debug|monitor_ready~q ),
	.take_action_ocimem_a(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|take_action_ocimem_a~1_combout ),
	.jdo_34(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[34]~q ),
	.writedata_0(\writedata[0]~q ),
	.take_action_ocireg(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|take_action_ocireg~0_combout ),
	.jdo_25(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[25]~q ),
	.jdo_21(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[20]~q ),
	.take_action_ocimem_a1(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|take_action_ocimem_a~combout ),
	.writedata_1(\writedata[1]~q ),
	.monitor_error1(\the_processor_nios2_gen2_0_cpu_nios2_oci_debug|monitor_error~q ),
	.jdo_19(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[18]~q ),
	.monitor_go1(\the_processor_nios2_gen2_0_cpu_nios2_oci_debug|monitor_go~q ),
	.jdo_23(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[23]~q ),
	.resetlatch1(\the_processor_nios2_gen2_0_cpu_nios2_oci_debug|resetlatch~q ),
	.jdo_24(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[24]~q ),
	.state_1(state_1),
	.clk_clk(clk_clk));

processor_processor_nios2_gen2_0_cpu_debug_slave_wrapper the_processor_nios2_gen2_0_cpu_debug_slave_wrapper(
	.sr_0(sr_0),
	.MonDReg_0(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[0]~q ),
	.MonDReg_4(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[4]~q ),
	.MonDReg_29(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[29]~q ),
	.MonDReg_5(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[5]~q ),
	.MonDReg_15(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[15]~q ),
	.MonDReg_12(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[12]~q ),
	.MonDReg_8(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[8]~q ),
	.MonDReg_18(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[18]~q ),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.break_readreg_0(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[0]~q ),
	.break_readreg_1(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[1]~q ),
	.MonDReg_1(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[1]~q ),
	.jdo_0(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[0]~q ),
	.jdo_36(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[36]~q ),
	.jdo_37(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[37]~q ),
	.ir_0(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|ir[0]~q ),
	.ir_1(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|ir[1]~q ),
	.enable_action_strobe(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|enable_action_strobe~q ),
	.jdo_3(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[3]~q ),
	.jdo_35(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[35]~q ),
	.take_action_ocimem_b(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|take_action_ocimem_b~combout ),
	.take_action_ocimem_a(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|take_action_ocimem_a~0_combout ),
	.monitor_ready(\the_processor_nios2_gen2_0_cpu_nios2_oci_debug|monitor_ready~q ),
	.hbreak_enabled(hbreak_enabled),
	.jdo_17(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[17]~q ),
	.take_action_ocimem_a1(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|take_action_ocimem_a~1_combout ),
	.jdo_34(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[34]~q ),
	.break_readreg_2(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[2]~q ),
	.MonDReg_2(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[2]~q ),
	.jdo_1(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[1]~q ),
	.jdo_4(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[4]~q ),
	.jdo_26(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[26]~q ),
	.jdo_28(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[28]~q ),
	.jdo_27(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[27]~q ),
	.jdo_25(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[25]~q ),
	.jdo_21(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[20]~q ),
	.take_action_ocimem_a2(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|take_action_ocimem_a~combout ),
	.jdo_33(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[33]~q ),
	.jdo_32(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[32]~q ),
	.jdo_31(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[31]~q ),
	.jdo_30(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[30]~q ),
	.jdo_29(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[29]~q ),
	.break_readreg_3(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[3]~q ),
	.MonDReg_3(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[3]~q ),
	.jdo_2(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[2]~q ),
	.jdo_5(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[5]~q ),
	.monitor_error(\the_processor_nios2_gen2_0_cpu_nios2_oci_debug|monitor_error~q ),
	.jdo_19(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[18]~q ),
	.break_readreg_16(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[16]~q ),
	.MonDReg_16(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[16]~q ),
	.break_readreg_4(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[4]~q ),
	.jdo_6(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[6]~q ),
	.break_readreg_25(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[25]~q ),
	.MonDReg_25(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[25]~q ),
	.break_readreg_27(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[27]~q ),
	.MonDReg_27(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[27]~q ),
	.break_readreg_26(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[26]~q ),
	.MonDReg_26(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[26]~q ),
	.break_readreg_24(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[24]~q ),
	.MonDReg_24(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[24]~q ),
	.break_readreg_20(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[20]~q ),
	.MonDReg_20(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[20]~q ),
	.break_readreg_19(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[19]~q ),
	.MonDReg_19(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[19]~q ),
	.MonDReg_22(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[22]~q ),
	.MonDReg_23(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[23]~q ),
	.jdo_23(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[23]~q ),
	.break_readreg_17(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[17]~q ),
	.MonDReg_17(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[17]~q ),
	.jdo_16(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[16]~q ),
	.resetlatch(\the_processor_nios2_gen2_0_cpu_nios2_oci_debug|resetlatch~q ),
	.break_readreg_31(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[31]~q ),
	.MonDReg_31(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[31]~q ),
	.break_readreg_30(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[30]~q ),
	.MonDReg_30(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[30]~q ),
	.break_readreg_29(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[29]~q ),
	.break_readreg_28(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[28]~q ),
	.MonDReg_28(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[28]~q ),
	.MonDReg_14(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[14]~q ),
	.MonDReg_11(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[11]~q ),
	.MonDReg_13(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[13]~q ),
	.MonDReg_10(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[10]~q ),
	.MonDReg_9(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[9]~q ),
	.MonDReg_7(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[7]~q ),
	.MonDReg_6(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[6]~q ),
	.MonDReg_21(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[21]~q ),
	.break_readreg_5(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[5]~q ),
	.jdo_7(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[7]~q ),
	.jdo_24(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[24]~q ),
	.break_readreg_18(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[18]~q ),
	.break_readreg_21(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[21]~q ),
	.jdo_22(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[22]~q ),
	.jdo_8(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[8]~q ),
	.jdo_14(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[14]~q ),
	.jdo_15(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[15]~q ),
	.jdo_13(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[13]~q ),
	.jdo_12(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[12]~q ),
	.jdo_11(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[11]~q ),
	.jdo_10(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[10]~q ),
	.jdo_9(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[9]~q ),
	.break_readreg_6(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[6]~q ),
	.break_readreg_22(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[22]~q ),
	.break_readreg_15(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[15]~q ),
	.break_readreg_7(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[7]~q ),
	.break_readreg_23(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[23]~q ),
	.break_readreg_13(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[13]~q ),
	.break_readreg_14(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[14]~q ),
	.break_readreg_12(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[12]~q ),
	.break_readreg_11(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[11]~q ),
	.break_readreg_10(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[10]~q ),
	.break_readreg_9(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[9]~q ),
	.break_readreg_8(\the_processor_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[8]~q ),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2),
	.clk_clk(clk_clk));

processor_processor_nios2_gen2_0_cpu_nios2_ocimem the_processor_nios2_gen2_0_cpu_nios2_ocimem(
	.MonDReg_0(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[0]~q ),
	.q_a_0(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ),
	.q_a_1(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ),
	.q_a_2(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ),
	.q_a_22(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_23(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_24(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ),
	.q_a_25(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ),
	.q_a_26(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ),
	.q_a_4(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ),
	.q_a_3(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ),
	.q_a_5(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_14(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_15(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_11(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_13(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_16(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ),
	.q_a_12(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_10(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_9(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_8(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_7(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ),
	.q_a_6(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ),
	.q_a_21(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ),
	.q_a_20(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ),
	.q_a_19(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ),
	.q_a_18(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ),
	.q_a_17(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ),
	.MonDReg_4(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[4]~q ),
	.MonDReg_29(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[29]~q ),
	.MonDReg_5(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[5]~q ),
	.MonDReg_15(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[15]~q ),
	.MonDReg_12(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[12]~q ),
	.q_a_27(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ),
	.q_a_28(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ),
	.q_a_29(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ),
	.q_a_30(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ),
	.q_a_31(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ),
	.MonDReg_8(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[8]~q ),
	.MonDReg_18(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[18]~q ),
	.waitrequest1(waitrequest),
	.write(\write~q ),
	.address_8(\address[8]~q ),
	.read(\read~q ),
	.MonDReg_1(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[1]~q ),
	.jdo_3(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[3]~q ),
	.jdo_35(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[35]~q ),
	.take_action_ocimem_b(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|take_action_ocimem_b~combout ),
	.take_action_ocimem_a(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|take_action_ocimem_a~0_combout ),
	.jdo_17(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[17]~q ),
	.take_action_ocimem_a1(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|take_action_ocimem_a~1_combout ),
	.jdo_34(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[34]~q ),
	.MonDReg_2(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[2]~q ),
	.jdo_4(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[4]~q ),
	.jdo_26(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[26]~q ),
	.jdo_28(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[28]~q ),
	.jdo_27(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[27]~q ),
	.debugaccess(\debugaccess~q ),
	.r_early_rst(r_early_rst),
	.writedata_0(\writedata[0]~q ),
	.address_0(\address[0]~q ),
	.address_1(\address[1]~q ),
	.address_2(\address[2]~q ),
	.address_3(\address[3]~q ),
	.address_4(\address[4]~q ),
	.address_5(\address[5]~q ),
	.address_6(\address[6]~q ),
	.address_7(\address[7]~q ),
	.byteenable_0(\byteenable[0]~q ),
	.jdo_25(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[25]~q ),
	.jdo_21(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[20]~q ),
	.jdo_33(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[33]~q ),
	.jdo_32(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[32]~q ),
	.jdo_31(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[31]~q ),
	.jdo_30(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[30]~q ),
	.jdo_29(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[29]~q ),
	.MonDReg_3(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[3]~q ),
	.jdo_5(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[5]~q ),
	.writedata_1(\writedata[1]~q ),
	.jdo_19(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[18]~q ),
	.writedata_3(\writedata[3]~q ),
	.MonDReg_16(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[16]~q ),
	.jdo_6(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[6]~q ),
	.writedata_2(\writedata[2]~q ),
	.MonDReg_25(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[25]~q ),
	.MonDReg_27(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[27]~q ),
	.MonDReg_26(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[26]~q ),
	.MonDReg_24(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[24]~q ),
	.MonDReg_20(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[20]~q ),
	.MonDReg_19(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[19]~q ),
	.MonDReg_22(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[22]~q ),
	.writedata_22(\writedata[22]~q ),
	.byteenable_2(\byteenable[2]~q ),
	.MonDReg_23(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[23]~q ),
	.writedata_23(\writedata[23]~q ),
	.writedata_24(\writedata[24]~q ),
	.byteenable_3(\byteenable[3]~q ),
	.writedata_25(\writedata[25]~q ),
	.writedata_26(\writedata[26]~q ),
	.writedata_4(\writedata[4]~q ),
	.jdo_23(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[23]~q ),
	.MonDReg_17(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[17]~q ),
	.jdo_16(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[16]~q ),
	.MonDReg_31(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[31]~q ),
	.MonDReg_30(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[30]~q ),
	.MonDReg_28(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[28]~q ),
	.writedata_5(\writedata[5]~q ),
	.MonDReg_14(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[14]~q ),
	.writedata_14(\writedata[14]~q ),
	.byteenable_1(\byteenable[1]~q ),
	.writedata_15(\writedata[15]~q ),
	.MonDReg_11(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[11]~q ),
	.writedata_11(\writedata[11]~q ),
	.MonDReg_13(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[13]~q ),
	.writedata_13(\writedata[13]~q ),
	.writedata_16(\writedata[16]~q ),
	.writedata_12(\writedata[12]~q ),
	.MonDReg_10(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[10]~q ),
	.writedata_10(\writedata[10]~q ),
	.MonDReg_9(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[9]~q ),
	.writedata_9(\writedata[9]~q ),
	.writedata_8(\writedata[8]~q ),
	.MonDReg_7(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[7]~q ),
	.writedata_7(\writedata[7]~q ),
	.MonDReg_6(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[6]~q ),
	.writedata_6(\writedata[6]~q ),
	.MonDReg_21(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[21]~q ),
	.writedata_21(\writedata[21]~q ),
	.writedata_20(\writedata[20]~q ),
	.writedata_19(\writedata[19]~q ),
	.writedata_18(\writedata[18]~q ),
	.writedata_17(\writedata[17]~q ),
	.jdo_7(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[7]~q ),
	.jdo_24(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[24]~q ),
	.jdo_22(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[22]~q ),
	.jdo_8(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[8]~q ),
	.jdo_14(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[14]~q ),
	.jdo_15(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[15]~q ),
	.writedata_27(\writedata[27]~q ),
	.writedata_28(\writedata[28]~q ),
	.writedata_29(\writedata[29]~q ),
	.writedata_30(\writedata[30]~q ),
	.writedata_31(\writedata[31]~q ),
	.jdo_13(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[13]~q ),
	.jdo_12(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[12]~q ),
	.jdo_11(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[11]~q ),
	.jdo_10(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[10]~q ),
	.jdo_9(\the_processor_nios2_gen2_0_cpu_debug_slave_wrapper|the_processor_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[9]~q ),
	.clk_clk(clk_clk));

processor_processor_nios2_gen2_0_cpu_nios2_avalon_reg the_processor_nios2_gen2_0_cpu_nios2_avalon_reg(
	.r_sync_rst(r_sync_rst),
	.write(\write~q ),
	.address_8(\address[8]~q ),
	.debugaccess(\debugaccess~q ),
	.writedata_0(\writedata[0]~q ),
	.address_0(\address[0]~q ),
	.address_1(\address[1]~q ),
	.address_2(\address[2]~q ),
	.address_3(\address[3]~q ),
	.address_4(\address[4]~q ),
	.address_5(\address[5]~q ),
	.address_6(\address[6]~q ),
	.address_7(\address[7]~q ),
	.Equal0(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal0~2_combout ),
	.take_action_ocireg(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|take_action_ocireg~0_combout ),
	.oci_ienable_0(oci_ienable_0),
	.oci_ienable_1(oci_ienable_1),
	.oci_single_step_mode1(oci_single_step_mode),
	.writedata_1(\writedata[1]~q ),
	.Equal1(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.writedata_3(\writedata[3]~q ),
	.oci_ienable_31(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ),
	.clk_clk(clk_clk));

dffeas write(
	.clk(clk_clk),
	.d(\write~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write~q ),
	.prn(vcc));
defparam write.is_wysiwyg = "true";
defparam write.power_up = "low";

dffeas read(
	.clk(clk_clk),
	.d(\read~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read~q ),
	.prn(vcc));
defparam read.is_wysiwyg = "true";
defparam read.power_up = "low";

cyclone10lp_lcell_comb \write~0 (
	.dataa(uav_write),
	.datab(saved_grant_0),
	.datac(mem_used_1),
	.datad(\write~q ),
	.cin(gnd),
	.combout(\write~0_combout ),
	.cout());
defparam \write~0 .lut_mask = 16'hEFFF;
defparam \write~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \write~1 (
	.dataa(waitrequest),
	.datab(WideOr1),
	.datac(\write~0_combout ),
	.datad(\write~q ),
	.cin(gnd),
	.combout(\write~1_combout ),
	.cout());
defparam \write~1 .lut_mask = 16'hFFFE;
defparam \write~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \read~0 (
	.dataa(waitrequest),
	.datab(\read~q ),
	.datac(rf_source_valid),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\read~0_combout ),
	.cout());
defparam \read~0 .lut_mask = 16'hB8FF;
defparam \read~0 .sum_lutc_input = "datac";

dffeas debugaccess(
	.clk(clk_clk),
	.d(debugaccess_nxt),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\debugaccess~q ),
	.prn(vcc));
defparam debugaccess.is_wysiwyg = "true";
defparam debugaccess.power_up = "low";

dffeas \writedata[0] (
	.clk(clk_clk),
	.d(writedata_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[0]~q ),
	.prn(vcc));
defparam \writedata[0] .is_wysiwyg = "true";
defparam \writedata[0] .power_up = "low";

dffeas \address[0] (
	.clk(clk_clk),
	.d(address_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[0]~q ),
	.prn(vcc));
defparam \address[0] .is_wysiwyg = "true";
defparam \address[0] .power_up = "low";

dffeas \address[1] (
	.clk(clk_clk),
	.d(address_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[1]~q ),
	.prn(vcc));
defparam \address[1] .is_wysiwyg = "true";
defparam \address[1] .power_up = "low";

dffeas \address[2] (
	.clk(clk_clk),
	.d(address_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[2]~q ),
	.prn(vcc));
defparam \address[2] .is_wysiwyg = "true";
defparam \address[2] .power_up = "low";

dffeas \address[3] (
	.clk(clk_clk),
	.d(address_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[3]~q ),
	.prn(vcc));
defparam \address[3] .is_wysiwyg = "true";
defparam \address[3] .power_up = "low";

dffeas \address[4] (
	.clk(clk_clk),
	.d(address_nxt[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[4]~q ),
	.prn(vcc));
defparam \address[4] .is_wysiwyg = "true";
defparam \address[4] .power_up = "low";

dffeas \address[5] (
	.clk(clk_clk),
	.d(address_nxt[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[5]~q ),
	.prn(vcc));
defparam \address[5] .is_wysiwyg = "true";
defparam \address[5] .power_up = "low";

dffeas \address[6] (
	.clk(clk_clk),
	.d(address_nxt[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[6]~q ),
	.prn(vcc));
defparam \address[6] .is_wysiwyg = "true";
defparam \address[6] .power_up = "low";

dffeas \address[7] (
	.clk(clk_clk),
	.d(address_nxt[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[7]~q ),
	.prn(vcc));
defparam \address[7] .is_wysiwyg = "true";
defparam \address[7] .power_up = "low";

dffeas \byteenable[0] (
	.clk(clk_clk),
	.d(byteenable_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[0]~q ),
	.prn(vcc));
defparam \byteenable[0] .is_wysiwyg = "true";
defparam \byteenable[0] .power_up = "low";

dffeas \writedata[1] (
	.clk(clk_clk),
	.d(writedata_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[1]~q ),
	.prn(vcc));
defparam \writedata[1] .is_wysiwyg = "true";
defparam \writedata[1] .power_up = "low";

dffeas \writedata[3] (
	.clk(clk_clk),
	.d(writedata_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[3]~q ),
	.prn(vcc));
defparam \writedata[3] .is_wysiwyg = "true";
defparam \writedata[3] .power_up = "low";

dffeas \writedata[2] (
	.clk(clk_clk),
	.d(writedata_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[2]~q ),
	.prn(vcc));
defparam \writedata[2] .is_wysiwyg = "true";
defparam \writedata[2] .power_up = "low";

dffeas \writedata[22] (
	.clk(clk_clk),
	.d(writedata_nxt[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[22]~q ),
	.prn(vcc));
defparam \writedata[22] .is_wysiwyg = "true";
defparam \writedata[22] .power_up = "low";

dffeas \byteenable[2] (
	.clk(clk_clk),
	.d(byteenable_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[2]~q ),
	.prn(vcc));
defparam \byteenable[2] .is_wysiwyg = "true";
defparam \byteenable[2] .power_up = "low";

dffeas \writedata[23] (
	.clk(clk_clk),
	.d(writedata_nxt[23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[23]~q ),
	.prn(vcc));
defparam \writedata[23] .is_wysiwyg = "true";
defparam \writedata[23] .power_up = "low";

dffeas \writedata[24] (
	.clk(clk_clk),
	.d(writedata_nxt[24]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[24]~q ),
	.prn(vcc));
defparam \writedata[24] .is_wysiwyg = "true";
defparam \writedata[24] .power_up = "low";

dffeas \byteenable[3] (
	.clk(clk_clk),
	.d(byteenable_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[3]~q ),
	.prn(vcc));
defparam \byteenable[3] .is_wysiwyg = "true";
defparam \byteenable[3] .power_up = "low";

dffeas \writedata[25] (
	.clk(clk_clk),
	.d(writedata_nxt[25]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[25]~q ),
	.prn(vcc));
defparam \writedata[25] .is_wysiwyg = "true";
defparam \writedata[25] .power_up = "low";

dffeas \writedata[26] (
	.clk(clk_clk),
	.d(writedata_nxt[26]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[26]~q ),
	.prn(vcc));
defparam \writedata[26] .is_wysiwyg = "true";
defparam \writedata[26] .power_up = "low";

dffeas \writedata[4] (
	.clk(clk_clk),
	.d(writedata_nxt[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[4]~q ),
	.prn(vcc));
defparam \writedata[4] .is_wysiwyg = "true";
defparam \writedata[4] .power_up = "low";

dffeas \writedata[5] (
	.clk(clk_clk),
	.d(writedata_nxt[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[5]~q ),
	.prn(vcc));
defparam \writedata[5] .is_wysiwyg = "true";
defparam \writedata[5] .power_up = "low";

dffeas \writedata[14] (
	.clk(clk_clk),
	.d(writedata_nxt[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[14]~q ),
	.prn(vcc));
defparam \writedata[14] .is_wysiwyg = "true";
defparam \writedata[14] .power_up = "low";

dffeas \byteenable[1] (
	.clk(clk_clk),
	.d(byteenable_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[1]~q ),
	.prn(vcc));
defparam \byteenable[1] .is_wysiwyg = "true";
defparam \byteenable[1] .power_up = "low";

dffeas \writedata[15] (
	.clk(clk_clk),
	.d(writedata_nxt[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[15]~q ),
	.prn(vcc));
defparam \writedata[15] .is_wysiwyg = "true";
defparam \writedata[15] .power_up = "low";

dffeas \writedata[11] (
	.clk(clk_clk),
	.d(writedata_nxt[11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[11]~q ),
	.prn(vcc));
defparam \writedata[11] .is_wysiwyg = "true";
defparam \writedata[11] .power_up = "low";

dffeas \writedata[13] (
	.clk(clk_clk),
	.d(writedata_nxt[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[13]~q ),
	.prn(vcc));
defparam \writedata[13] .is_wysiwyg = "true";
defparam \writedata[13] .power_up = "low";

dffeas \writedata[16] (
	.clk(clk_clk),
	.d(writedata_nxt[16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[16]~q ),
	.prn(vcc));
defparam \writedata[16] .is_wysiwyg = "true";
defparam \writedata[16] .power_up = "low";

dffeas \writedata[12] (
	.clk(clk_clk),
	.d(writedata_nxt[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[12]~q ),
	.prn(vcc));
defparam \writedata[12] .is_wysiwyg = "true";
defparam \writedata[12] .power_up = "low";

dffeas \writedata[10] (
	.clk(clk_clk),
	.d(writedata_nxt[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[10]~q ),
	.prn(vcc));
defparam \writedata[10] .is_wysiwyg = "true";
defparam \writedata[10] .power_up = "low";

dffeas \writedata[9] (
	.clk(clk_clk),
	.d(writedata_nxt[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[9]~q ),
	.prn(vcc));
defparam \writedata[9] .is_wysiwyg = "true";
defparam \writedata[9] .power_up = "low";

dffeas \writedata[8] (
	.clk(clk_clk),
	.d(writedata_nxt[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[8]~q ),
	.prn(vcc));
defparam \writedata[8] .is_wysiwyg = "true";
defparam \writedata[8] .power_up = "low";

dffeas \writedata[7] (
	.clk(clk_clk),
	.d(writedata_nxt[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[7]~q ),
	.prn(vcc));
defparam \writedata[7] .is_wysiwyg = "true";
defparam \writedata[7] .power_up = "low";

dffeas \writedata[6] (
	.clk(clk_clk),
	.d(writedata_nxt[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[6]~q ),
	.prn(vcc));
defparam \writedata[6] .is_wysiwyg = "true";
defparam \writedata[6] .power_up = "low";

dffeas \writedata[21] (
	.clk(clk_clk),
	.d(writedata_nxt[21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[21]~q ),
	.prn(vcc));
defparam \writedata[21] .is_wysiwyg = "true";
defparam \writedata[21] .power_up = "low";

dffeas \writedata[20] (
	.clk(clk_clk),
	.d(writedata_nxt[20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[20]~q ),
	.prn(vcc));
defparam \writedata[20] .is_wysiwyg = "true";
defparam \writedata[20] .power_up = "low";

dffeas \writedata[19] (
	.clk(clk_clk),
	.d(writedata_nxt[19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[19]~q ),
	.prn(vcc));
defparam \writedata[19] .is_wysiwyg = "true";
defparam \writedata[19] .power_up = "low";

dffeas \writedata[18] (
	.clk(clk_clk),
	.d(writedata_nxt[18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[18]~q ),
	.prn(vcc));
defparam \writedata[18] .is_wysiwyg = "true";
defparam \writedata[18] .power_up = "low";

dffeas \writedata[17] (
	.clk(clk_clk),
	.d(writedata_nxt[17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[17]~q ),
	.prn(vcc));
defparam \writedata[17] .is_wysiwyg = "true";
defparam \writedata[17] .power_up = "low";

dffeas \writedata[27] (
	.clk(clk_clk),
	.d(writedata_nxt[27]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[27]~q ),
	.prn(vcc));
defparam \writedata[27] .is_wysiwyg = "true";
defparam \writedata[27] .power_up = "low";

dffeas \writedata[28] (
	.clk(clk_clk),
	.d(writedata_nxt[28]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[28]~q ),
	.prn(vcc));
defparam \writedata[28] .is_wysiwyg = "true";
defparam \writedata[28] .power_up = "low";

dffeas \writedata[29] (
	.clk(clk_clk),
	.d(writedata_nxt[29]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[29]~q ),
	.prn(vcc));
defparam \writedata[29] .is_wysiwyg = "true";
defparam \writedata[29] .power_up = "low";

dffeas \writedata[30] (
	.clk(clk_clk),
	.d(writedata_nxt[30]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[30]~q ),
	.prn(vcc));
defparam \writedata[30] .is_wysiwyg = "true";
defparam \writedata[30] .power_up = "low";

dffeas \writedata[31] (
	.clk(clk_clk),
	.d(writedata_nxt[31]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[31]~q ),
	.prn(vcc));
defparam \writedata[31] .is_wysiwyg = "true";
defparam \writedata[31] .power_up = "low";

dffeas \readdata[0] (
	.clk(clk_clk),
	.d(\readdata~0_combout ),
	.asdata(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk_clk),
	.d(\readdata~6_combout ),
	.asdata(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk_clk),
	.d(\readdata~8_combout ),
	.asdata(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk_clk),
	.d(\readdata~9_combout ),
	.asdata(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[22] (
	.clk(clk_clk),
	.d(\readdata~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_22),
	.prn(vcc));
defparam \readdata[22] .is_wysiwyg = "true";
defparam \readdata[22] .power_up = "low";

dffeas \readdata[23] (
	.clk(clk_clk),
	.d(\readdata~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_23),
	.prn(vcc));
defparam \readdata[23] .is_wysiwyg = "true";
defparam \readdata[23] .power_up = "low";

dffeas \readdata[24] (
	.clk(clk_clk),
	.d(\readdata~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_24),
	.prn(vcc));
defparam \readdata[24] .is_wysiwyg = "true";
defparam \readdata[24] .power_up = "low";

dffeas \readdata[25] (
	.clk(clk_clk),
	.d(\readdata~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_25),
	.prn(vcc));
defparam \readdata[25] .is_wysiwyg = "true";
defparam \readdata[25] .power_up = "low";

dffeas \readdata[26] (
	.clk(clk_clk),
	.d(\readdata~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_26),
	.prn(vcc));
defparam \readdata[26] .is_wysiwyg = "true";
defparam \readdata[26] .power_up = "low";

dffeas \readdata[4] (
	.clk(clk_clk),
	.d(\readdata~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[5] (
	.clk(clk_clk),
	.d(\readdata~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[14] (
	.clk(clk_clk),
	.d(\readdata~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_14),
	.prn(vcc));
defparam \readdata[14] .is_wysiwyg = "true";
defparam \readdata[14] .power_up = "low";

dffeas \readdata[15] (
	.clk(clk_clk),
	.d(\readdata~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_15),
	.prn(vcc));
defparam \readdata[15] .is_wysiwyg = "true";
defparam \readdata[15] .power_up = "low";

dffeas \readdata[11] (
	.clk(clk_clk),
	.d(\readdata~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_11),
	.prn(vcc));
defparam \readdata[11] .is_wysiwyg = "true";
defparam \readdata[11] .power_up = "low";

dffeas \readdata[13] (
	.clk(clk_clk),
	.d(\readdata~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_13),
	.prn(vcc));
defparam \readdata[13] .is_wysiwyg = "true";
defparam \readdata[13] .power_up = "low";

dffeas \readdata[16] (
	.clk(clk_clk),
	.d(\readdata~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_16),
	.prn(vcc));
defparam \readdata[16] .is_wysiwyg = "true";
defparam \readdata[16] .power_up = "low";

dffeas \readdata[12] (
	.clk(clk_clk),
	.d(\readdata~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_12),
	.prn(vcc));
defparam \readdata[12] .is_wysiwyg = "true";
defparam \readdata[12] .power_up = "low";

dffeas \readdata[10] (
	.clk(clk_clk),
	.d(\readdata~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_10),
	.prn(vcc));
defparam \readdata[10] .is_wysiwyg = "true";
defparam \readdata[10] .power_up = "low";

dffeas \readdata[9] (
	.clk(clk_clk),
	.d(\readdata~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_9),
	.prn(vcc));
defparam \readdata[9] .is_wysiwyg = "true";
defparam \readdata[9] .power_up = "low";

dffeas \readdata[8] (
	.clk(clk_clk),
	.d(\readdata~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_8),
	.prn(vcc));
defparam \readdata[8] .is_wysiwyg = "true";
defparam \readdata[8] .power_up = "low";

dffeas \readdata[7] (
	.clk(clk_clk),
	.d(\readdata~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_7),
	.prn(vcc));
defparam \readdata[7] .is_wysiwyg = "true";
defparam \readdata[7] .power_up = "low";

dffeas \readdata[6] (
	.clk(clk_clk),
	.d(\readdata~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

dffeas \readdata[21] (
	.clk(clk_clk),
	.d(\readdata~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_21),
	.prn(vcc));
defparam \readdata[21] .is_wysiwyg = "true";
defparam \readdata[21] .power_up = "low";

dffeas \readdata[20] (
	.clk(clk_clk),
	.d(\readdata~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_20),
	.prn(vcc));
defparam \readdata[20] .is_wysiwyg = "true";
defparam \readdata[20] .power_up = "low";

dffeas \readdata[19] (
	.clk(clk_clk),
	.d(\readdata~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_19),
	.prn(vcc));
defparam \readdata[19] .is_wysiwyg = "true";
defparam \readdata[19] .power_up = "low";

dffeas \readdata[18] (
	.clk(clk_clk),
	.d(\readdata~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_18),
	.prn(vcc));
defparam \readdata[18] .is_wysiwyg = "true";
defparam \readdata[18] .power_up = "low";

dffeas \readdata[17] (
	.clk(clk_clk),
	.d(\readdata~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_17),
	.prn(vcc));
defparam \readdata[17] .is_wysiwyg = "true";
defparam \readdata[17] .power_up = "low";

dffeas \readdata[27] (
	.clk(clk_clk),
	.d(\readdata~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_27),
	.prn(vcc));
defparam \readdata[27] .is_wysiwyg = "true";
defparam \readdata[27] .power_up = "low";

dffeas \readdata[28] (
	.clk(clk_clk),
	.d(\readdata~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_28),
	.prn(vcc));
defparam \readdata[28] .is_wysiwyg = "true";
defparam \readdata[28] .power_up = "low";

dffeas \readdata[29] (
	.clk(clk_clk),
	.d(\readdata~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_29),
	.prn(vcc));
defparam \readdata[29] .is_wysiwyg = "true";
defparam \readdata[29] .power_up = "low";

dffeas \readdata[30] (
	.clk(clk_clk),
	.d(\readdata~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_30),
	.prn(vcc));
defparam \readdata[30] .is_wysiwyg = "true";
defparam \readdata[30] .power_up = "low";

dffeas \readdata[31] (
	.clk(clk_clk),
	.d(\readdata~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_31),
	.prn(vcc));
defparam \readdata[31] .is_wysiwyg = "true";
defparam \readdata[31] .power_up = "low";

cyclone10lp_lcell_comb \readdata~0 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_oci_debug|monitor_error~q ),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal0~2_combout ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datad(oci_ienable_0),
	.cin(gnd),
	.combout(\readdata~0_combout ),
	.cout());
defparam \readdata~0 .lut_mask = 16'hB8FF;
defparam \readdata~0 .sum_lutc_input = "datac";

dffeas \address[8] (
	.clk(clk_clk),
	.d(address_nxt[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[8]~q ),
	.prn(vcc));
defparam \address[8] .is_wysiwyg = "true";
defparam \address[8] .power_up = "low";

cyclone10lp_lcell_comb \readdata~6 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_oci_debug|monitor_ready~q ),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal0~2_combout ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datad(oci_ienable_1),
	.cin(gnd),
	.combout(\readdata~6_combout ),
	.cout());
defparam \readdata~6 .lut_mask = 16'hB8FF;
defparam \readdata~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata~8 (
	.dataa(oci_single_step_mode),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ),
	.datad(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal0~2_combout ),
	.cin(gnd),
	.combout(\readdata~8_combout ),
	.cout());
defparam \readdata~8 .lut_mask = 16'hFAFC;
defparam \readdata~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata~9 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_oci_debug|monitor_go~q ),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ),
	.datad(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal0~2_combout ),
	.cin(gnd),
	.combout(\readdata~9_combout ),
	.cout());
defparam \readdata~9 .lut_mask = 16'hFAFC;
defparam \readdata~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata~1 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~1_combout ),
	.cout());
defparam \readdata~1 .lut_mask = 16'hFAFC;
defparam \readdata~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata~2 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~2_combout ),
	.cout());
defparam \readdata~2 .lut_mask = 16'hFAFC;
defparam \readdata~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata~3 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~3_combout ),
	.cout());
defparam \readdata~3 .lut_mask = 16'hFAFC;
defparam \readdata~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata~4 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~4_combout ),
	.cout());
defparam \readdata~4 .lut_mask = 16'hFAFC;
defparam \readdata~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata~5 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~5_combout ),
	.cout());
defparam \readdata~5 .lut_mask = 16'hFAFC;
defparam \readdata~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata~7 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~7_combout ),
	.cout());
defparam \readdata~7 .lut_mask = 16'hFAFC;
defparam \readdata~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata~10 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~10_combout ),
	.cout());
defparam \readdata~10 .lut_mask = 16'hFAFC;
defparam \readdata~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata~11 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~11_combout ),
	.cout());
defparam \readdata~11 .lut_mask = 16'hFAFC;
defparam \readdata~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata~12 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~12_combout ),
	.cout());
defparam \readdata~12 .lut_mask = 16'hFAFC;
defparam \readdata~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata~13 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~13_combout ),
	.cout());
defparam \readdata~13 .lut_mask = 16'hFAFC;
defparam \readdata~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata~14 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~14_combout ),
	.cout());
defparam \readdata~14 .lut_mask = 16'hFAFC;
defparam \readdata~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata~15 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~15_combout ),
	.cout());
defparam \readdata~15 .lut_mask = 16'hFAFC;
defparam \readdata~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata~16 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~16_combout ),
	.cout());
defparam \readdata~16 .lut_mask = 16'hFAFC;
defparam \readdata~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata~17 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~17_combout ),
	.cout());
defparam \readdata~17 .lut_mask = 16'hFAFC;
defparam \readdata~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata~18 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~18_combout ),
	.cout());
defparam \readdata~18 .lut_mask = 16'hFAFC;
defparam \readdata~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata~19 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~19_combout ),
	.cout());
defparam \readdata~19 .lut_mask = 16'hFAFC;
defparam \readdata~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata~20 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~20_combout ),
	.cout());
defparam \readdata~20 .lut_mask = 16'hFAFC;
defparam \readdata~20 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata~21 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~21_combout ),
	.cout());
defparam \readdata~21 .lut_mask = 16'hFAFC;
defparam \readdata~21 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata~22 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~22_combout ),
	.cout());
defparam \readdata~22 .lut_mask = 16'hFAFC;
defparam \readdata~22 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata~23 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~23_combout ),
	.cout());
defparam \readdata~23 .lut_mask = 16'hFAFC;
defparam \readdata~23 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata~24 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~24_combout ),
	.cout());
defparam \readdata~24 .lut_mask = 16'hFAFC;
defparam \readdata~24 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata~25 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~25_combout ),
	.cout());
defparam \readdata~25 .lut_mask = 16'hFAFC;
defparam \readdata~25 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata~26 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~26_combout ),
	.cout());
defparam \readdata~26 .lut_mask = 16'hFAFC;
defparam \readdata~26 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata~27 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~27_combout ),
	.cout());
defparam \readdata~27 .lut_mask = 16'hFAFC;
defparam \readdata~27 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata~28 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~28_combout ),
	.cout());
defparam \readdata~28 .lut_mask = 16'hFAFC;
defparam \readdata~28 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata~29 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~29_combout ),
	.cout());
defparam \readdata~29 .lut_mask = 16'hFAFC;
defparam \readdata~29 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata~30 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~30_combout ),
	.cout());
defparam \readdata~30 .lut_mask = 16'hFAFC;
defparam \readdata~30 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata~31 (
	.dataa(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_processor_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[31]~q ),
	.datac(\the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~31_combout ),
	.cout());
defparam \readdata~31 .lut_mask = 16'hFAFC;
defparam \readdata~31 .sum_lutc_input = "datac";

endmodule

module processor_processor_nios2_gen2_0_cpu_debug_slave_wrapper (
	sr_0,
	MonDReg_0,
	MonDReg_4,
	MonDReg_29,
	MonDReg_5,
	MonDReg_15,
	MonDReg_12,
	MonDReg_8,
	MonDReg_18,
	ir_out_0,
	ir_out_1,
	break_readreg_0,
	break_readreg_1,
	MonDReg_1,
	jdo_0,
	jdo_36,
	jdo_37,
	ir_0,
	ir_1,
	enable_action_strobe,
	jdo_3,
	jdo_35,
	take_action_ocimem_b,
	take_action_ocimem_a,
	monitor_ready,
	hbreak_enabled,
	jdo_17,
	take_action_ocimem_a1,
	jdo_34,
	break_readreg_2,
	MonDReg_2,
	jdo_1,
	jdo_4,
	jdo_26,
	jdo_28,
	jdo_27,
	jdo_25,
	jdo_21,
	jdo_20,
	take_action_ocimem_a2,
	jdo_33,
	jdo_32,
	jdo_31,
	jdo_30,
	jdo_29,
	break_readreg_3,
	MonDReg_3,
	jdo_2,
	jdo_5,
	monitor_error,
	jdo_19,
	jdo_18,
	break_readreg_16,
	MonDReg_16,
	break_readreg_4,
	jdo_6,
	break_readreg_25,
	MonDReg_25,
	break_readreg_27,
	MonDReg_27,
	break_readreg_26,
	MonDReg_26,
	break_readreg_24,
	MonDReg_24,
	break_readreg_20,
	MonDReg_20,
	break_readreg_19,
	MonDReg_19,
	MonDReg_22,
	MonDReg_23,
	jdo_23,
	break_readreg_17,
	MonDReg_17,
	jdo_16,
	resetlatch,
	break_readreg_31,
	MonDReg_31,
	break_readreg_30,
	MonDReg_30,
	break_readreg_29,
	break_readreg_28,
	MonDReg_28,
	MonDReg_14,
	MonDReg_11,
	MonDReg_13,
	MonDReg_10,
	MonDReg_9,
	MonDReg_7,
	MonDReg_6,
	MonDReg_21,
	break_readreg_5,
	jdo_7,
	jdo_24,
	break_readreg_18,
	break_readreg_21,
	jdo_22,
	jdo_8,
	jdo_14,
	jdo_15,
	jdo_13,
	jdo_12,
	jdo_11,
	jdo_10,
	jdo_9,
	break_readreg_6,
	break_readreg_22,
	break_readreg_15,
	break_readreg_7,
	break_readreg_23,
	break_readreg_13,
	break_readreg_14,
	break_readreg_12,
	break_readreg_11,
	break_readreg_10,
	break_readreg_9,
	break_readreg_8,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	sr_0;
input 	MonDReg_0;
input 	MonDReg_4;
input 	MonDReg_29;
input 	MonDReg_5;
input 	MonDReg_15;
input 	MonDReg_12;
input 	MonDReg_8;
input 	MonDReg_18;
output 	ir_out_0;
output 	ir_out_1;
input 	break_readreg_0;
input 	break_readreg_1;
input 	MonDReg_1;
output 	jdo_0;
output 	jdo_36;
output 	jdo_37;
output 	ir_0;
output 	ir_1;
output 	enable_action_strobe;
output 	jdo_3;
output 	jdo_35;
output 	take_action_ocimem_b;
output 	take_action_ocimem_a;
input 	monitor_ready;
input 	hbreak_enabled;
output 	jdo_17;
output 	take_action_ocimem_a1;
output 	jdo_34;
input 	break_readreg_2;
input 	MonDReg_2;
output 	jdo_1;
output 	jdo_4;
output 	jdo_26;
output 	jdo_28;
output 	jdo_27;
output 	jdo_25;
output 	jdo_21;
output 	jdo_20;
output 	take_action_ocimem_a2;
output 	jdo_33;
output 	jdo_32;
output 	jdo_31;
output 	jdo_30;
output 	jdo_29;
input 	break_readreg_3;
input 	MonDReg_3;
output 	jdo_2;
output 	jdo_5;
input 	monitor_error;
output 	jdo_19;
output 	jdo_18;
input 	break_readreg_16;
input 	MonDReg_16;
input 	break_readreg_4;
output 	jdo_6;
input 	break_readreg_25;
input 	MonDReg_25;
input 	break_readreg_27;
input 	MonDReg_27;
input 	break_readreg_26;
input 	MonDReg_26;
input 	break_readreg_24;
input 	MonDReg_24;
input 	break_readreg_20;
input 	MonDReg_20;
input 	break_readreg_19;
input 	MonDReg_19;
input 	MonDReg_22;
input 	MonDReg_23;
output 	jdo_23;
input 	break_readreg_17;
input 	MonDReg_17;
output 	jdo_16;
input 	resetlatch;
input 	break_readreg_31;
input 	MonDReg_31;
input 	break_readreg_30;
input 	MonDReg_30;
input 	break_readreg_29;
input 	break_readreg_28;
input 	MonDReg_28;
input 	MonDReg_14;
input 	MonDReg_11;
input 	MonDReg_13;
input 	MonDReg_10;
input 	MonDReg_9;
input 	MonDReg_7;
input 	MonDReg_6;
input 	MonDReg_21;
input 	break_readreg_5;
output 	jdo_7;
output 	jdo_24;
input 	break_readreg_18;
input 	break_readreg_21;
output 	jdo_22;
output 	jdo_8;
output 	jdo_14;
output 	jdo_15;
output 	jdo_13;
output 	jdo_12;
output 	jdo_11;
output 	jdo_10;
output 	jdo_9;
input 	break_readreg_6;
input 	break_readreg_22;
input 	break_readreg_15;
input 	break_readreg_7;
input 	break_readreg_23;
input 	break_readreg_13;
input 	break_readreg_14;
input 	break_readreg_12;
input 	break_readreg_11;
input 	break_readreg_10;
input 	break_readreg_9;
input 	break_readreg_8;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[35]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[31]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[7]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[15]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[1]~q ;
wire \processor_nios2_gen2_0_cpu_debug_slave_phy|virtual_state_cdr~combout ;
wire \processor_nios2_gen2_0_cpu_debug_slave_phy|virtual_state_sdr~0_combout ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[2]~q ;
wire \processor_nios2_gen2_0_cpu_debug_slave_phy|virtual_state_uir~0_combout ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[3]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[4]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[36]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[37]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[17]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[34]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[5]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[26]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[28]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[27]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[25]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[21]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[20]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[18]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[33]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[32]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[30]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[29]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[6]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[19]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[22]~q ;
wire \processor_nios2_gen2_0_cpu_debug_slave_phy|virtual_state_udr~0_combout ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[23]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[16]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[8]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[24]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[14]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[13]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[12]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[11]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[10]~q ;
wire \the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[9]~q ;


processor_sld_virtual_jtag_basic_1 processor_nios2_gen2_0_cpu_debug_slave_phy(
	.virtual_state_cdr1(\processor_nios2_gen2_0_cpu_debug_slave_phy|virtual_state_cdr~combout ),
	.virtual_state_sdr(\processor_nios2_gen2_0_cpu_debug_slave_phy|virtual_state_sdr~0_combout ),
	.virtual_state_uir(\processor_nios2_gen2_0_cpu_debug_slave_phy|virtual_state_uir~0_combout ),
	.virtual_state_udr(\processor_nios2_gen2_0_cpu_debug_slave_phy|virtual_state_udr~0_combout ),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3));

processor_processor_nios2_gen2_0_cpu_debug_slave_sysclk the_processor_nios2_gen2_0_cpu_debug_slave_sysclk(
	.sr_0(sr_0),
	.sr_35(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[35]~q ),
	.sr_31(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[31]~q ),
	.sr_7(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[7]~q ),
	.sr_15(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[15]~q ),
	.sr_1(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[1]~q ),
	.sr_2(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[2]~q ),
	.virtual_state_uir(\processor_nios2_gen2_0_cpu_debug_slave_phy|virtual_state_uir~0_combout ),
	.sr_3(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[3]~q ),
	.jdo_0(jdo_0),
	.jdo_36(jdo_36),
	.jdo_37(jdo_37),
	.ir_0(ir_0),
	.ir_1(ir_1),
	.enable_action_strobe1(enable_action_strobe),
	.jdo_3(jdo_3),
	.jdo_35(jdo_35),
	.take_action_ocimem_b1(take_action_ocimem_b),
	.take_action_ocimem_a1(take_action_ocimem_a),
	.jdo_17(jdo_17),
	.take_action_ocimem_a2(take_action_ocimem_a1),
	.jdo_34(jdo_34),
	.sr_4(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[4]~q ),
	.jdo_1(jdo_1),
	.jdo_4(jdo_4),
	.sr_36(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[36]~q ),
	.sr_37(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[37]~q ),
	.jdo_26(jdo_26),
	.jdo_28(jdo_28),
	.jdo_27(jdo_27),
	.jdo_25(jdo_25),
	.jdo_21(jdo_21),
	.jdo_20(jdo_20),
	.take_action_ocimem_a3(take_action_ocimem_a2),
	.sr_17(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[17]~q ),
	.jdo_33(jdo_33),
	.jdo_32(jdo_32),
	.jdo_31(jdo_31),
	.jdo_30(jdo_30),
	.jdo_29(jdo_29),
	.sr_34(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[34]~q ),
	.sr_5(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[5]~q ),
	.jdo_2(jdo_2),
	.jdo_5(jdo_5),
	.sr_26(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[26]~q ),
	.sr_28(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[28]~q ),
	.sr_27(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[27]~q ),
	.sr_25(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[25]~q ),
	.jdo_19(jdo_19),
	.jdo_18(jdo_18),
	.sr_21(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[21]~q ),
	.sr_20(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[20]~q ),
	.sr_18(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[18]~q ),
	.sr_33(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[33]~q ),
	.sr_32(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[32]~q ),
	.sr_30(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[30]~q ),
	.sr_29(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[29]~q ),
	.sr_6(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[6]~q ),
	.jdo_6(jdo_6),
	.sr_19(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[19]~q ),
	.sr_22(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[22]~q ),
	.jdo_23(jdo_23),
	.jdo_16(jdo_16),
	.jdo_7(jdo_7),
	.virtual_state_udr(\processor_nios2_gen2_0_cpu_debug_slave_phy|virtual_state_udr~0_combout ),
	.jdo_24(jdo_24),
	.sr_23(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[23]~q ),
	.jdo_22(jdo_22),
	.sr_16(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[16]~q ),
	.jdo_8(jdo_8),
	.jdo_14(jdo_14),
	.jdo_15(jdo_15),
	.jdo_13(jdo_13),
	.jdo_12(jdo_12),
	.jdo_11(jdo_11),
	.jdo_10(jdo_10),
	.jdo_9(jdo_9),
	.sr_8(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[8]~q ),
	.sr_24(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[24]~q ),
	.sr_14(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[14]~q ),
	.sr_13(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[13]~q ),
	.sr_12(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[12]~q ),
	.sr_11(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[11]~q ),
	.sr_10(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[10]~q ),
	.sr_9(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[9]~q ),
	.ir_in({irf_reg_1_2,irf_reg_0_2}),
	.clk_clk(clk_clk));

processor_processor_nios2_gen2_0_cpu_debug_slave_tck the_processor_nios2_gen2_0_cpu_debug_slave_tck(
	.sr_0(sr_0),
	.MonDReg_0(MonDReg_0),
	.sr_35(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[35]~q ),
	.sr_31(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[31]~q ),
	.MonDReg_4(MonDReg_4),
	.MonDReg_29(MonDReg_29),
	.MonDReg_5(MonDReg_5),
	.MonDReg_15(MonDReg_15),
	.MonDReg_12(MonDReg_12),
	.MonDReg_8(MonDReg_8),
	.MonDReg_18(MonDReg_18),
	.sr_7(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[7]~q ),
	.sr_15(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[15]~q ),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.sr_1(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[1]~q ),
	.virtual_state_cdr(\processor_nios2_gen2_0_cpu_debug_slave_phy|virtual_state_cdr~combout ),
	.virtual_state_sdr(\processor_nios2_gen2_0_cpu_debug_slave_phy|virtual_state_sdr~0_combout ),
	.sr_2(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[2]~q ),
	.break_readreg_0(break_readreg_0),
	.virtual_state_uir(\processor_nios2_gen2_0_cpu_debug_slave_phy|virtual_state_uir~0_combout ),
	.sr_3(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[3]~q ),
	.break_readreg_1(break_readreg_1),
	.MonDReg_1(MonDReg_1),
	.monitor_ready(monitor_ready),
	.hbreak_enabled(hbreak_enabled),
	.sr_4(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[4]~q ),
	.break_readreg_2(break_readreg_2),
	.MonDReg_2(MonDReg_2),
	.sr_36(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[36]~q ),
	.sr_37(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[37]~q ),
	.sr_17(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[17]~q ),
	.sr_34(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[34]~q ),
	.sr_5(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[5]~q ),
	.break_readreg_3(break_readreg_3),
	.MonDReg_3(MonDReg_3),
	.sr_26(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[26]~q ),
	.sr_28(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[28]~q ),
	.sr_27(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[27]~q ),
	.sr_25(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[25]~q ),
	.monitor_error(monitor_error),
	.sr_21(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[21]~q ),
	.sr_20(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[20]~q ),
	.sr_18(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[18]~q ),
	.break_readreg_16(break_readreg_16),
	.MonDReg_16(MonDReg_16),
	.sr_33(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[33]~q ),
	.sr_32(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[32]~q ),
	.sr_30(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[30]~q ),
	.sr_29(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[29]~q ),
	.sr_6(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[6]~q ),
	.break_readreg_4(break_readreg_4),
	.break_readreg_25(break_readreg_25),
	.MonDReg_25(MonDReg_25),
	.break_readreg_27(break_readreg_27),
	.MonDReg_27(MonDReg_27),
	.break_readreg_26(break_readreg_26),
	.MonDReg_26(MonDReg_26),
	.break_readreg_24(break_readreg_24),
	.MonDReg_24(MonDReg_24),
	.sr_19(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[19]~q ),
	.sr_22(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[22]~q ),
	.break_readreg_20(break_readreg_20),
	.MonDReg_20(MonDReg_20),
	.break_readreg_19(break_readreg_19),
	.MonDReg_19(MonDReg_19),
	.MonDReg_22(MonDReg_22),
	.MonDReg_23(MonDReg_23),
	.break_readreg_17(break_readreg_17),
	.MonDReg_17(MonDReg_17),
	.resetlatch(resetlatch),
	.break_readreg_31(break_readreg_31),
	.MonDReg_31(MonDReg_31),
	.break_readreg_30(break_readreg_30),
	.MonDReg_30(MonDReg_30),
	.break_readreg_29(break_readreg_29),
	.break_readreg_28(break_readreg_28),
	.MonDReg_28(MonDReg_28),
	.MonDReg_14(MonDReg_14),
	.MonDReg_11(MonDReg_11),
	.MonDReg_13(MonDReg_13),
	.MonDReg_10(MonDReg_10),
	.MonDReg_9(MonDReg_9),
	.MonDReg_7(MonDReg_7),
	.MonDReg_6(MonDReg_6),
	.MonDReg_21(MonDReg_21),
	.break_readreg_5(break_readreg_5),
	.break_readreg_18(break_readreg_18),
	.sr_23(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[23]~q ),
	.break_readreg_21(break_readreg_21),
	.sr_16(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[16]~q ),
	.break_readreg_6(break_readreg_6),
	.sr_8(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[8]~q ),
	.sr_24(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[24]~q ),
	.break_readreg_22(break_readreg_22),
	.break_readreg_15(break_readreg_15),
	.sr_14(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[14]~q ),
	.sr_13(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[13]~q ),
	.sr_12(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[12]~q ),
	.sr_11(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[11]~q ),
	.sr_10(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[10]~q ),
	.sr_9(\the_processor_nios2_gen2_0_cpu_debug_slave_tck|sr[9]~q ),
	.break_readreg_7(break_readreg_7),
	.break_readreg_23(break_readreg_23),
	.break_readreg_13(break_readreg_13),
	.break_readreg_14(break_readreg_14),
	.break_readreg_12(break_readreg_12),
	.break_readreg_11(break_readreg_11),
	.break_readreg_10(break_readreg_10),
	.break_readreg_9(break_readreg_9),
	.break_readreg_8(break_readreg_8),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2));

endmodule

module processor_processor_nios2_gen2_0_cpu_debug_slave_sysclk (
	sr_0,
	sr_35,
	sr_31,
	sr_7,
	sr_15,
	sr_1,
	sr_2,
	virtual_state_uir,
	sr_3,
	jdo_0,
	jdo_36,
	jdo_37,
	ir_0,
	ir_1,
	enable_action_strobe1,
	jdo_3,
	jdo_35,
	take_action_ocimem_b1,
	take_action_ocimem_a1,
	jdo_17,
	take_action_ocimem_a2,
	jdo_34,
	sr_4,
	jdo_1,
	jdo_4,
	sr_36,
	sr_37,
	jdo_26,
	jdo_28,
	jdo_27,
	jdo_25,
	jdo_21,
	jdo_20,
	take_action_ocimem_a3,
	sr_17,
	jdo_33,
	jdo_32,
	jdo_31,
	jdo_30,
	jdo_29,
	sr_34,
	sr_5,
	jdo_2,
	jdo_5,
	sr_26,
	sr_28,
	sr_27,
	sr_25,
	jdo_19,
	jdo_18,
	sr_21,
	sr_20,
	sr_18,
	sr_33,
	sr_32,
	sr_30,
	sr_29,
	sr_6,
	jdo_6,
	sr_19,
	sr_22,
	jdo_23,
	jdo_16,
	jdo_7,
	virtual_state_udr,
	jdo_24,
	sr_23,
	jdo_22,
	sr_16,
	jdo_8,
	jdo_14,
	jdo_15,
	jdo_13,
	jdo_12,
	jdo_11,
	jdo_10,
	jdo_9,
	sr_8,
	sr_24,
	sr_14,
	sr_13,
	sr_12,
	sr_11,
	sr_10,
	sr_9,
	ir_in,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	sr_0;
input 	sr_35;
input 	sr_31;
input 	sr_7;
input 	sr_15;
input 	sr_1;
input 	sr_2;
input 	virtual_state_uir;
input 	sr_3;
output 	jdo_0;
output 	jdo_36;
output 	jdo_37;
output 	ir_0;
output 	ir_1;
output 	enable_action_strobe1;
output 	jdo_3;
output 	jdo_35;
output 	take_action_ocimem_b1;
output 	take_action_ocimem_a1;
output 	jdo_17;
output 	take_action_ocimem_a2;
output 	jdo_34;
input 	sr_4;
output 	jdo_1;
output 	jdo_4;
input 	sr_36;
input 	sr_37;
output 	jdo_26;
output 	jdo_28;
output 	jdo_27;
output 	jdo_25;
output 	jdo_21;
output 	jdo_20;
output 	take_action_ocimem_a3;
input 	sr_17;
output 	jdo_33;
output 	jdo_32;
output 	jdo_31;
output 	jdo_30;
output 	jdo_29;
input 	sr_34;
input 	sr_5;
output 	jdo_2;
output 	jdo_5;
input 	sr_26;
input 	sr_28;
input 	sr_27;
input 	sr_25;
output 	jdo_19;
output 	jdo_18;
input 	sr_21;
input 	sr_20;
input 	sr_18;
input 	sr_33;
input 	sr_32;
input 	sr_30;
input 	sr_29;
input 	sr_6;
output 	jdo_6;
input 	sr_19;
input 	sr_22;
output 	jdo_23;
output 	jdo_16;
output 	jdo_7;
input 	virtual_state_udr;
output 	jdo_24;
input 	sr_23;
output 	jdo_22;
input 	sr_16;
output 	jdo_8;
output 	jdo_14;
output 	jdo_15;
output 	jdo_13;
output 	jdo_12;
output 	jdo_11;
output 	jdo_10;
output 	jdo_9;
input 	sr_8;
input 	sr_24;
input 	sr_14;
input 	sr_13;
input 	sr_12;
input 	sr_11;
input 	sr_10;
input 	sr_9;
input 	[1:0] ir_in;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer3|dreg[0]~q ;
wire \the_altera_std_synchronizer4|dreg[0]~q ;
wire \sync2_udr~q ;
wire \update_jdo_strobe~0_combout ;
wire \update_jdo_strobe~q ;
wire \sync2_uir~q ;
wire \jxuir~0_combout ;
wire \jxuir~q ;


processor_altera_std_synchronizer_1 the_altera_std_synchronizer4(
	.din(virtual_state_uir),
	.dreg_0(\the_altera_std_synchronizer4|dreg[0]~q ),
	.clk(clk_clk));

processor_altera_std_synchronizer the_altera_std_synchronizer3(
	.dreg_0(\the_altera_std_synchronizer3|dreg[0]~q ),
	.din(virtual_state_udr),
	.clk(clk_clk));

dffeas \jdo[0] (
	.clk(clk_clk),
	.d(sr_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_0),
	.prn(vcc));
defparam \jdo[0] .is_wysiwyg = "true";
defparam \jdo[0] .power_up = "low";

dffeas \jdo[36] (
	.clk(clk_clk),
	.d(sr_36),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_36),
	.prn(vcc));
defparam \jdo[36] .is_wysiwyg = "true";
defparam \jdo[36] .power_up = "low";

dffeas \jdo[37] (
	.clk(clk_clk),
	.d(sr_37),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_37),
	.prn(vcc));
defparam \jdo[37] .is_wysiwyg = "true";
defparam \jdo[37] .power_up = "low";

dffeas \ir[0] (
	.clk(clk_clk),
	.d(ir_in[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\jxuir~q ),
	.q(ir_0),
	.prn(vcc));
defparam \ir[0] .is_wysiwyg = "true";
defparam \ir[0] .power_up = "low";

dffeas \ir[1] (
	.clk(clk_clk),
	.d(ir_in[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\jxuir~q ),
	.q(ir_1),
	.prn(vcc));
defparam \ir[1] .is_wysiwyg = "true";
defparam \ir[1] .power_up = "low";

dffeas enable_action_strobe(
	.clk(clk_clk),
	.d(\update_jdo_strobe~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(enable_action_strobe1),
	.prn(vcc));
defparam enable_action_strobe.is_wysiwyg = "true";
defparam enable_action_strobe.power_up = "low";

dffeas \jdo[3] (
	.clk(clk_clk),
	.d(sr_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_3),
	.prn(vcc));
defparam \jdo[3] .is_wysiwyg = "true";
defparam \jdo[3] .power_up = "low";

dffeas \jdo[35] (
	.clk(clk_clk),
	.d(sr_35),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_35),
	.prn(vcc));
defparam \jdo[35] .is_wysiwyg = "true";
defparam \jdo[35] .power_up = "low";

cyclone10lp_lcell_comb take_action_ocimem_b(
	.dataa(enable_action_strobe1),
	.datab(jdo_35),
	.datac(ir_1),
	.datad(ir_0),
	.cin(gnd),
	.combout(take_action_ocimem_b1),
	.cout());
defparam take_action_ocimem_b.lut_mask = 16'hEFFF;
defparam take_action_ocimem_b.sum_lutc_input = "datac";

cyclone10lp_lcell_comb \take_action_ocimem_a~0 (
	.dataa(enable_action_strobe1),
	.datab(gnd),
	.datac(ir_1),
	.datad(ir_0),
	.cin(gnd),
	.combout(take_action_ocimem_a1),
	.cout());
defparam \take_action_ocimem_a~0 .lut_mask = 16'hAFFF;
defparam \take_action_ocimem_a~0 .sum_lutc_input = "datac";

dffeas \jdo[17] (
	.clk(clk_clk),
	.d(sr_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_17),
	.prn(vcc));
defparam \jdo[17] .is_wysiwyg = "true";
defparam \jdo[17] .power_up = "low";

cyclone10lp_lcell_comb \take_action_ocimem_a~1 (
	.dataa(enable_action_strobe1),
	.datab(ir_1),
	.datac(ir_0),
	.datad(jdo_35),
	.cin(gnd),
	.combout(take_action_ocimem_a2),
	.cout());
defparam \take_action_ocimem_a~1 .lut_mask = 16'hBFFF;
defparam \take_action_ocimem_a~1 .sum_lutc_input = "datac";

dffeas \jdo[34] (
	.clk(clk_clk),
	.d(sr_34),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_34),
	.prn(vcc));
defparam \jdo[34] .is_wysiwyg = "true";
defparam \jdo[34] .power_up = "low";

dffeas \jdo[1] (
	.clk(clk_clk),
	.d(sr_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_1),
	.prn(vcc));
defparam \jdo[1] .is_wysiwyg = "true";
defparam \jdo[1] .power_up = "low";

dffeas \jdo[4] (
	.clk(clk_clk),
	.d(sr_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_4),
	.prn(vcc));
defparam \jdo[4] .is_wysiwyg = "true";
defparam \jdo[4] .power_up = "low";

dffeas \jdo[26] (
	.clk(clk_clk),
	.d(sr_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_26),
	.prn(vcc));
defparam \jdo[26] .is_wysiwyg = "true";
defparam \jdo[26] .power_up = "low";

dffeas \jdo[28] (
	.clk(clk_clk),
	.d(sr_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_28),
	.prn(vcc));
defparam \jdo[28] .is_wysiwyg = "true";
defparam \jdo[28] .power_up = "low";

dffeas \jdo[27] (
	.clk(clk_clk),
	.d(sr_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_27),
	.prn(vcc));
defparam \jdo[27] .is_wysiwyg = "true";
defparam \jdo[27] .power_up = "low";

dffeas \jdo[25] (
	.clk(clk_clk),
	.d(sr_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_25),
	.prn(vcc));
defparam \jdo[25] .is_wysiwyg = "true";
defparam \jdo[25] .power_up = "low";

dffeas \jdo[21] (
	.clk(clk_clk),
	.d(sr_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_21),
	.prn(vcc));
defparam \jdo[21] .is_wysiwyg = "true";
defparam \jdo[21] .power_up = "low";

dffeas \jdo[20] (
	.clk(clk_clk),
	.d(sr_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_20),
	.prn(vcc));
defparam \jdo[20] .is_wysiwyg = "true";
defparam \jdo[20] .power_up = "low";

cyclone10lp_lcell_comb take_action_ocimem_a(
	.dataa(take_action_ocimem_a1),
	.datab(jdo_34),
	.datac(gnd),
	.datad(jdo_35),
	.cin(gnd),
	.combout(take_action_ocimem_a3),
	.cout());
defparam take_action_ocimem_a.lut_mask = 16'hEEFF;
defparam take_action_ocimem_a.sum_lutc_input = "datac";

dffeas \jdo[33] (
	.clk(clk_clk),
	.d(sr_33),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_33),
	.prn(vcc));
defparam \jdo[33] .is_wysiwyg = "true";
defparam \jdo[33] .power_up = "low";

dffeas \jdo[32] (
	.clk(clk_clk),
	.d(sr_32),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_32),
	.prn(vcc));
defparam \jdo[32] .is_wysiwyg = "true";
defparam \jdo[32] .power_up = "low";

dffeas \jdo[31] (
	.clk(clk_clk),
	.d(sr_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_31),
	.prn(vcc));
defparam \jdo[31] .is_wysiwyg = "true";
defparam \jdo[31] .power_up = "low";

dffeas \jdo[30] (
	.clk(clk_clk),
	.d(sr_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_30),
	.prn(vcc));
defparam \jdo[30] .is_wysiwyg = "true";
defparam \jdo[30] .power_up = "low";

dffeas \jdo[29] (
	.clk(clk_clk),
	.d(sr_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_29),
	.prn(vcc));
defparam \jdo[29] .is_wysiwyg = "true";
defparam \jdo[29] .power_up = "low";

dffeas \jdo[2] (
	.clk(clk_clk),
	.d(sr_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_2),
	.prn(vcc));
defparam \jdo[2] .is_wysiwyg = "true";
defparam \jdo[2] .power_up = "low";

dffeas \jdo[5] (
	.clk(clk_clk),
	.d(sr_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_5),
	.prn(vcc));
defparam \jdo[5] .is_wysiwyg = "true";
defparam \jdo[5] .power_up = "low";

dffeas \jdo[19] (
	.clk(clk_clk),
	.d(sr_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_19),
	.prn(vcc));
defparam \jdo[19] .is_wysiwyg = "true";
defparam \jdo[19] .power_up = "low";

dffeas \jdo[18] (
	.clk(clk_clk),
	.d(sr_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_18),
	.prn(vcc));
defparam \jdo[18] .is_wysiwyg = "true";
defparam \jdo[18] .power_up = "low";

dffeas \jdo[6] (
	.clk(clk_clk),
	.d(sr_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_6),
	.prn(vcc));
defparam \jdo[6] .is_wysiwyg = "true";
defparam \jdo[6] .power_up = "low";

dffeas \jdo[23] (
	.clk(clk_clk),
	.d(sr_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_23),
	.prn(vcc));
defparam \jdo[23] .is_wysiwyg = "true";
defparam \jdo[23] .power_up = "low";

dffeas \jdo[16] (
	.clk(clk_clk),
	.d(sr_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_16),
	.prn(vcc));
defparam \jdo[16] .is_wysiwyg = "true";
defparam \jdo[16] .power_up = "low";

dffeas \jdo[7] (
	.clk(clk_clk),
	.d(sr_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_7),
	.prn(vcc));
defparam \jdo[7] .is_wysiwyg = "true";
defparam \jdo[7] .power_up = "low";

dffeas \jdo[24] (
	.clk(clk_clk),
	.d(sr_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_24),
	.prn(vcc));
defparam \jdo[24] .is_wysiwyg = "true";
defparam \jdo[24] .power_up = "low";

dffeas \jdo[22] (
	.clk(clk_clk),
	.d(sr_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_22),
	.prn(vcc));
defparam \jdo[22] .is_wysiwyg = "true";
defparam \jdo[22] .power_up = "low";

dffeas \jdo[8] (
	.clk(clk_clk),
	.d(sr_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_8),
	.prn(vcc));
defparam \jdo[8] .is_wysiwyg = "true";
defparam \jdo[8] .power_up = "low";

dffeas \jdo[14] (
	.clk(clk_clk),
	.d(sr_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_14),
	.prn(vcc));
defparam \jdo[14] .is_wysiwyg = "true";
defparam \jdo[14] .power_up = "low";

dffeas \jdo[15] (
	.clk(clk_clk),
	.d(sr_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_15),
	.prn(vcc));
defparam \jdo[15] .is_wysiwyg = "true";
defparam \jdo[15] .power_up = "low";

dffeas \jdo[13] (
	.clk(clk_clk),
	.d(sr_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_13),
	.prn(vcc));
defparam \jdo[13] .is_wysiwyg = "true";
defparam \jdo[13] .power_up = "low";

dffeas \jdo[12] (
	.clk(clk_clk),
	.d(sr_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_12),
	.prn(vcc));
defparam \jdo[12] .is_wysiwyg = "true";
defparam \jdo[12] .power_up = "low";

dffeas \jdo[11] (
	.clk(clk_clk),
	.d(sr_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_11),
	.prn(vcc));
defparam \jdo[11] .is_wysiwyg = "true";
defparam \jdo[11] .power_up = "low";

dffeas \jdo[10] (
	.clk(clk_clk),
	.d(sr_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_10),
	.prn(vcc));
defparam \jdo[10] .is_wysiwyg = "true";
defparam \jdo[10] .power_up = "low";

dffeas \jdo[9] (
	.clk(clk_clk),
	.d(sr_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_9),
	.prn(vcc));
defparam \jdo[9] .is_wysiwyg = "true";
defparam \jdo[9] .power_up = "low";

dffeas sync2_udr(
	.clk(clk_clk),
	.d(\the_altera_std_synchronizer3|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sync2_udr~q ),
	.prn(vcc));
defparam sync2_udr.is_wysiwyg = "true";
defparam sync2_udr.power_up = "low";

cyclone10lp_lcell_comb \update_jdo_strobe~0 (
	.dataa(\the_altera_std_synchronizer3|dreg[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\sync2_udr~q ),
	.cin(gnd),
	.combout(\update_jdo_strobe~0_combout ),
	.cout());
defparam \update_jdo_strobe~0 .lut_mask = 16'hAAFF;
defparam \update_jdo_strobe~0 .sum_lutc_input = "datac";

dffeas update_jdo_strobe(
	.clk(clk_clk),
	.d(\update_jdo_strobe~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\update_jdo_strobe~q ),
	.prn(vcc));
defparam update_jdo_strobe.is_wysiwyg = "true";
defparam update_jdo_strobe.power_up = "low";

dffeas sync2_uir(
	.clk(clk_clk),
	.d(\the_altera_std_synchronizer4|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sync2_uir~q ),
	.prn(vcc));
defparam sync2_uir.is_wysiwyg = "true";
defparam sync2_uir.power_up = "low";

cyclone10lp_lcell_comb \jxuir~0 (
	.dataa(\the_altera_std_synchronizer4|dreg[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\sync2_uir~q ),
	.cin(gnd),
	.combout(\jxuir~0_combout ),
	.cout());
defparam \jxuir~0 .lut_mask = 16'hAAFF;
defparam \jxuir~0 .sum_lutc_input = "datac";

dffeas jxuir(
	.clk(clk_clk),
	.d(\jxuir~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jxuir~q ),
	.prn(vcc));
defparam jxuir.is_wysiwyg = "true";
defparam jxuir.power_up = "low";

endmodule

module processor_altera_std_synchronizer (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module processor_altera_std_synchronizer_1 (
	din,
	dreg_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	din;
output 	dreg_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module processor_processor_nios2_gen2_0_cpu_debug_slave_tck (
	sr_0,
	MonDReg_0,
	sr_35,
	sr_31,
	MonDReg_4,
	MonDReg_29,
	MonDReg_5,
	MonDReg_15,
	MonDReg_12,
	MonDReg_8,
	MonDReg_18,
	sr_7,
	sr_15,
	ir_out_0,
	ir_out_1,
	sr_1,
	virtual_state_cdr,
	virtual_state_sdr,
	sr_2,
	break_readreg_0,
	virtual_state_uir,
	sr_3,
	break_readreg_1,
	MonDReg_1,
	monitor_ready,
	hbreak_enabled,
	sr_4,
	break_readreg_2,
	MonDReg_2,
	sr_36,
	sr_37,
	sr_17,
	sr_34,
	sr_5,
	break_readreg_3,
	MonDReg_3,
	sr_26,
	sr_28,
	sr_27,
	sr_25,
	monitor_error,
	sr_21,
	sr_20,
	sr_18,
	break_readreg_16,
	MonDReg_16,
	sr_33,
	sr_32,
	sr_30,
	sr_29,
	sr_6,
	break_readreg_4,
	break_readreg_25,
	MonDReg_25,
	break_readreg_27,
	MonDReg_27,
	break_readreg_26,
	MonDReg_26,
	break_readreg_24,
	MonDReg_24,
	sr_19,
	sr_22,
	break_readreg_20,
	MonDReg_20,
	break_readreg_19,
	MonDReg_19,
	MonDReg_22,
	MonDReg_23,
	break_readreg_17,
	MonDReg_17,
	resetlatch,
	break_readreg_31,
	MonDReg_31,
	break_readreg_30,
	MonDReg_30,
	break_readreg_29,
	break_readreg_28,
	MonDReg_28,
	MonDReg_14,
	MonDReg_11,
	MonDReg_13,
	MonDReg_10,
	MonDReg_9,
	MonDReg_7,
	MonDReg_6,
	MonDReg_21,
	break_readreg_5,
	break_readreg_18,
	sr_23,
	break_readreg_21,
	sr_16,
	break_readreg_6,
	sr_8,
	sr_24,
	break_readreg_22,
	break_readreg_15,
	sr_14,
	sr_13,
	sr_12,
	sr_11,
	sr_10,
	sr_9,
	break_readreg_7,
	break_readreg_23,
	break_readreg_13,
	break_readreg_14,
	break_readreg_12,
	break_readreg_11,
	break_readreg_10,
	break_readreg_9,
	break_readreg_8,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2)/* synthesis synthesis_greybox=1 */;
output 	sr_0;
input 	MonDReg_0;
output 	sr_35;
output 	sr_31;
input 	MonDReg_4;
input 	MonDReg_29;
input 	MonDReg_5;
input 	MonDReg_15;
input 	MonDReg_12;
input 	MonDReg_8;
input 	MonDReg_18;
output 	sr_7;
output 	sr_15;
output 	ir_out_0;
output 	ir_out_1;
output 	sr_1;
input 	virtual_state_cdr;
input 	virtual_state_sdr;
output 	sr_2;
input 	break_readreg_0;
input 	virtual_state_uir;
output 	sr_3;
input 	break_readreg_1;
input 	MonDReg_1;
input 	monitor_ready;
input 	hbreak_enabled;
output 	sr_4;
input 	break_readreg_2;
input 	MonDReg_2;
output 	sr_36;
output 	sr_37;
output 	sr_17;
output 	sr_34;
output 	sr_5;
input 	break_readreg_3;
input 	MonDReg_3;
output 	sr_26;
output 	sr_28;
output 	sr_27;
output 	sr_25;
input 	monitor_error;
output 	sr_21;
output 	sr_20;
output 	sr_18;
input 	break_readreg_16;
input 	MonDReg_16;
output 	sr_33;
output 	sr_32;
output 	sr_30;
output 	sr_29;
output 	sr_6;
input 	break_readreg_4;
input 	break_readreg_25;
input 	MonDReg_25;
input 	break_readreg_27;
input 	MonDReg_27;
input 	break_readreg_26;
input 	MonDReg_26;
input 	break_readreg_24;
input 	MonDReg_24;
output 	sr_19;
output 	sr_22;
input 	break_readreg_20;
input 	MonDReg_20;
input 	break_readreg_19;
input 	MonDReg_19;
input 	MonDReg_22;
input 	MonDReg_23;
input 	break_readreg_17;
input 	MonDReg_17;
input 	resetlatch;
input 	break_readreg_31;
input 	MonDReg_31;
input 	break_readreg_30;
input 	MonDReg_30;
input 	break_readreg_29;
input 	break_readreg_28;
input 	MonDReg_28;
input 	MonDReg_14;
input 	MonDReg_11;
input 	MonDReg_13;
input 	MonDReg_10;
input 	MonDReg_9;
input 	MonDReg_7;
input 	MonDReg_6;
input 	MonDReg_21;
input 	break_readreg_5;
input 	break_readreg_18;
output 	sr_23;
input 	break_readreg_21;
output 	sr_16;
input 	break_readreg_6;
output 	sr_8;
output 	sr_24;
input 	break_readreg_22;
input 	break_readreg_15;
output 	sr_14;
output 	sr_13;
output 	sr_12;
output 	sr_11;
output 	sr_10;
output 	sr_9;
input 	break_readreg_7;
input 	break_readreg_23;
input 	break_readreg_13;
input 	break_readreg_14;
input 	break_readreg_12;
input 	break_readreg_11;
input 	break_readreg_10;
input 	break_readreg_9;
input 	break_readreg_8;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer2|dreg[0]~q ;
wire \the_altera_std_synchronizer1|dreg[0]~q ;
wire \DRsize.000~q ;
wire \sr[0]~5_combout ;
wire \Mux37~0_combout ;
wire \sr~10_combout ;
wire \DRsize.100~q ;
wire \sr[35]~6_combout ;
wire \sr~23_combout ;
wire \sr~24_combout ;
wire \sr~25_combout ;
wire \sr[31]~50_combout ;
wire \sr[31]~7_combout ;
wire \Mux30~0_combout ;
wire \sr[7]~8_combout ;
wire \sr[33]~83_combout ;
wire \DRsize.010~q ;
wire \sr[15]~9_combout ;
wire \sr~71_combout ;
wire \sr~72_combout ;
wire \sr~11_combout ;
wire \sr~12_combout ;
wire \sr[13]~13_combout ;
wire \sr~14_combout ;
wire \sr~15_combout ;
wire \sr~16_combout ;
wire \sr~17_combout ;
wire \sr~18_combout ;
wire \sr~19_combout ;
wire \sr~20_combout ;
wire \sr[36]~21_combout ;
wire \sr~22_combout ;
wire \sr~26_combout ;
wire \sr~27_combout ;
wire \sr~28_combout ;
wire \sr[33]~29_combout ;
wire \sr~30_combout ;
wire \sr~31_combout ;
wire \sr~32_combout ;
wire \sr~33_combout ;
wire \sr~34_combout ;
wire \sr~35_combout ;
wire \sr~36_combout ;
wire \sr~37_combout ;
wire \sr~38_combout ;
wire \sr~39_combout ;
wire \sr~40_combout ;
wire \sr~41_combout ;
wire \sr~42_combout ;
wire \sr~43_combout ;
wire \sr~44_combout ;
wire \sr~45_combout ;
wire \sr~46_combout ;
wire \sr~47_combout ;
wire \sr~48_combout ;
wire \sr~49_combout ;
wire \sr~51_combout ;
wire \sr~52_combout ;
wire \sr~53_combout ;
wire \sr~54_combout ;
wire \sr~55_combout ;
wire \sr~56_combout ;
wire \sr~57_combout ;
wire \sr~58_combout ;
wire \sr~59_combout ;
wire \sr~60_combout ;
wire \sr~61_combout ;
wire \sr~62_combout ;
wire \sr~63_combout ;
wire \sr~64_combout ;
wire \sr~65_combout ;
wire \sr~66_combout ;
wire \sr~67_combout ;
wire \sr~68_combout ;
wire \sr~69_combout ;
wire \sr~70_combout ;
wire \sr~73_combout ;
wire \sr~74_combout ;
wire \sr~75_combout ;
wire \sr~76_combout ;
wire \sr~77_combout ;
wire \sr~78_combout ;
wire \sr~79_combout ;
wire \sr~80_combout ;
wire \sr~81_combout ;
wire \sr~82_combout ;


processor_altera_std_synchronizer_3 the_altera_std_synchronizer2(
	.dreg_0(\the_altera_std_synchronizer2|dreg[0]~q ),
	.din(monitor_ready),
	.clk(altera_internal_jtag));

processor_altera_std_synchronizer_2 the_altera_std_synchronizer1(
	.dreg_0(\the_altera_std_synchronizer1|dreg[0]~q ),
	.din(hbreak_enabled),
	.clk(altera_internal_jtag));

dffeas \sr[0] (
	.clk(altera_internal_jtag),
	.d(\sr[0]~5_combout ),
	.asdata(\sr~10_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!virtual_state_sdr),
	.ena(vcc),
	.q(sr_0),
	.prn(vcc));
defparam \sr[0] .is_wysiwyg = "true";
defparam \sr[0] .power_up = "low";

dffeas \sr[35] (
	.clk(altera_internal_jtag),
	.d(\sr[35]~6_combout ),
	.asdata(\sr~25_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!virtual_state_sdr),
	.ena(vcc),
	.q(sr_35),
	.prn(vcc));
defparam \sr[35] .is_wysiwyg = "true";
defparam \sr[35] .power_up = "low";

dffeas \sr[31] (
	.clk(altera_internal_jtag),
	.d(\sr[31]~7_combout ),
	.asdata(sr_32),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(virtual_state_sdr),
	.ena(vcc),
	.q(sr_31),
	.prn(vcc));
defparam \sr[31] .is_wysiwyg = "true";
defparam \sr[31] .power_up = "low";

dffeas \sr[7] (
	.clk(altera_internal_jtag),
	.d(\sr[7]~8_combout ),
	.asdata(sr_8),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(virtual_state_sdr),
	.ena(vcc),
	.q(sr_7),
	.prn(vcc));
defparam \sr[7] .is_wysiwyg = "true";
defparam \sr[7] .power_up = "low";

dffeas \sr[15] (
	.clk(altera_internal_jtag),
	.d(\sr[15]~9_combout ),
	.asdata(\sr~72_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!virtual_state_sdr),
	.ena(vcc),
	.q(sr_15),
	.prn(vcc));
defparam \sr[15] .is_wysiwyg = "true";
defparam \sr[15] .power_up = "low";

dffeas \ir_out[0] (
	.clk(altera_internal_jtag),
	.d(\the_altera_std_synchronizer2|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ir_out_0),
	.prn(vcc));
defparam \ir_out[0] .is_wysiwyg = "true";
defparam \ir_out[0] .power_up = "low";

dffeas \ir_out[1] (
	.clk(altera_internal_jtag),
	.d(\the_altera_std_synchronizer1|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ir_out_1),
	.prn(vcc));
defparam \ir_out[1] .is_wysiwyg = "true";
defparam \ir_out[1] .power_up = "low";

dffeas \sr[1] (
	.clk(altera_internal_jtag),
	.d(\sr~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[13]~13_combout ),
	.q(sr_1),
	.prn(vcc));
defparam \sr[1] .is_wysiwyg = "true";
defparam \sr[1] .power_up = "low";

dffeas \sr[2] (
	.clk(altera_internal_jtag),
	.d(\sr~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[13]~13_combout ),
	.q(sr_2),
	.prn(vcc));
defparam \sr[2] .is_wysiwyg = "true";
defparam \sr[2] .power_up = "low";

dffeas \sr[3] (
	.clk(altera_internal_jtag),
	.d(\sr~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[13]~13_combout ),
	.q(sr_3),
	.prn(vcc));
defparam \sr[3] .is_wysiwyg = "true";
defparam \sr[3] .power_up = "low";

dffeas \sr[4] (
	.clk(altera_internal_jtag),
	.d(\sr~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[13]~13_combout ),
	.q(sr_4),
	.prn(vcc));
defparam \sr[4] .is_wysiwyg = "true";
defparam \sr[4] .power_up = "low";

dffeas \sr[36] (
	.clk(altera_internal_jtag),
	.d(\sr~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[36]~21_combout ),
	.q(sr_36),
	.prn(vcc));
defparam \sr[36] .is_wysiwyg = "true";
defparam \sr[36] .power_up = "low";

dffeas \sr[37] (
	.clk(altera_internal_jtag),
	.d(\sr~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[36]~21_combout ),
	.q(sr_37),
	.prn(vcc));
defparam \sr[37] .is_wysiwyg = "true";
defparam \sr[37] .power_up = "low";

dffeas \sr[17] (
	.clk(altera_internal_jtag),
	.d(\sr~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_17),
	.prn(vcc));
defparam \sr[17] .is_wysiwyg = "true";
defparam \sr[17] .power_up = "low";

dffeas \sr[34] (
	.clk(altera_internal_jtag),
	.d(\sr~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_34),
	.prn(vcc));
defparam \sr[34] .is_wysiwyg = "true";
defparam \sr[34] .power_up = "low";

dffeas \sr[5] (
	.clk(altera_internal_jtag),
	.d(\sr~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[13]~13_combout ),
	.q(sr_5),
	.prn(vcc));
defparam \sr[5] .is_wysiwyg = "true";
defparam \sr[5] .power_up = "low";

dffeas \sr[26] (
	.clk(altera_internal_jtag),
	.d(\sr~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_26),
	.prn(vcc));
defparam \sr[26] .is_wysiwyg = "true";
defparam \sr[26] .power_up = "low";

dffeas \sr[28] (
	.clk(altera_internal_jtag),
	.d(\sr~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_28),
	.prn(vcc));
defparam \sr[28] .is_wysiwyg = "true";
defparam \sr[28] .power_up = "low";

dffeas \sr[27] (
	.clk(altera_internal_jtag),
	.d(\sr~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_27),
	.prn(vcc));
defparam \sr[27] .is_wysiwyg = "true";
defparam \sr[27] .power_up = "low";

dffeas \sr[25] (
	.clk(altera_internal_jtag),
	.d(\sr~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_25),
	.prn(vcc));
defparam \sr[25] .is_wysiwyg = "true";
defparam \sr[25] .power_up = "low";

dffeas \sr[21] (
	.clk(altera_internal_jtag),
	.d(\sr~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_21),
	.prn(vcc));
defparam \sr[21] .is_wysiwyg = "true";
defparam \sr[21] .power_up = "low";

dffeas \sr[20] (
	.clk(altera_internal_jtag),
	.d(\sr~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_20),
	.prn(vcc));
defparam \sr[20] .is_wysiwyg = "true";
defparam \sr[20] .power_up = "low";

dffeas \sr[18] (
	.clk(altera_internal_jtag),
	.d(\sr~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_18),
	.prn(vcc));
defparam \sr[18] .is_wysiwyg = "true";
defparam \sr[18] .power_up = "low";

dffeas \sr[33] (
	.clk(altera_internal_jtag),
	.d(\sr~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_33),
	.prn(vcc));
defparam \sr[33] .is_wysiwyg = "true";
defparam \sr[33] .power_up = "low";

dffeas \sr[32] (
	.clk(altera_internal_jtag),
	.d(\sr~49_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_32),
	.prn(vcc));
defparam \sr[32] .is_wysiwyg = "true";
defparam \sr[32] .power_up = "low";

dffeas \sr[30] (
	.clk(altera_internal_jtag),
	.d(\sr~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_30),
	.prn(vcc));
defparam \sr[30] .is_wysiwyg = "true";
defparam \sr[30] .power_up = "low";

dffeas \sr[29] (
	.clk(altera_internal_jtag),
	.d(\sr~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_29),
	.prn(vcc));
defparam \sr[29] .is_wysiwyg = "true";
defparam \sr[29] .power_up = "low";

dffeas \sr[6] (
	.clk(altera_internal_jtag),
	.d(\sr~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[13]~13_combout ),
	.q(sr_6),
	.prn(vcc));
defparam \sr[6] .is_wysiwyg = "true";
defparam \sr[6] .power_up = "low";

dffeas \sr[19] (
	.clk(altera_internal_jtag),
	.d(\sr~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_19),
	.prn(vcc));
defparam \sr[19] .is_wysiwyg = "true";
defparam \sr[19] .power_up = "low";

dffeas \sr[22] (
	.clk(altera_internal_jtag),
	.d(\sr~60_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_22),
	.prn(vcc));
defparam \sr[22] .is_wysiwyg = "true";
defparam \sr[22] .power_up = "low";

dffeas \sr[23] (
	.clk(altera_internal_jtag),
	.d(\sr~62_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_23),
	.prn(vcc));
defparam \sr[23] .is_wysiwyg = "true";
defparam \sr[23] .power_up = "low";

dffeas \sr[16] (
	.clk(altera_internal_jtag),
	.d(\sr~64_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_16),
	.prn(vcc));
defparam \sr[16] .is_wysiwyg = "true";
defparam \sr[16] .power_up = "low";

dffeas \sr[8] (
	.clk(altera_internal_jtag),
	.d(\sr~66_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[13]~13_combout ),
	.q(sr_8),
	.prn(vcc));
defparam \sr[8] .is_wysiwyg = "true";
defparam \sr[8] .power_up = "low";

dffeas \sr[24] (
	.clk(altera_internal_jtag),
	.d(\sr~68_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_24),
	.prn(vcc));
defparam \sr[24] .is_wysiwyg = "true";
defparam \sr[24] .power_up = "low";

dffeas \sr[14] (
	.clk(altera_internal_jtag),
	.d(\sr~70_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[13]~13_combout ),
	.q(sr_14),
	.prn(vcc));
defparam \sr[14] .is_wysiwyg = "true";
defparam \sr[14] .power_up = "low";

dffeas \sr[13] (
	.clk(altera_internal_jtag),
	.d(\sr~74_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[13]~13_combout ),
	.q(sr_13),
	.prn(vcc));
defparam \sr[13] .is_wysiwyg = "true";
defparam \sr[13] .power_up = "low";

dffeas \sr[12] (
	.clk(altera_internal_jtag),
	.d(\sr~76_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[13]~13_combout ),
	.q(sr_12),
	.prn(vcc));
defparam \sr[12] .is_wysiwyg = "true";
defparam \sr[12] .power_up = "low";

dffeas \sr[11] (
	.clk(altera_internal_jtag),
	.d(\sr~78_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[13]~13_combout ),
	.q(sr_11),
	.prn(vcc));
defparam \sr[11] .is_wysiwyg = "true";
defparam \sr[11] .power_up = "low";

dffeas \sr[10] (
	.clk(altera_internal_jtag),
	.d(\sr~80_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[13]~13_combout ),
	.q(sr_10),
	.prn(vcc));
defparam \sr[10] .is_wysiwyg = "true";
defparam \sr[10] .power_up = "low";

dffeas \sr[9] (
	.clk(altera_internal_jtag),
	.d(\sr~82_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[13]~13_combout ),
	.q(sr_9),
	.prn(vcc));
defparam \sr[9] .is_wysiwyg = "true";
defparam \sr[9] .power_up = "low";

dffeas \DRsize.000 (
	.clk(altera_internal_jtag),
	.d(vcc),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.000~q ),
	.prn(vcc));
defparam \DRsize.000 .is_wysiwyg = "true";
defparam \DRsize.000 .power_up = "low";

cyclone10lp_lcell_comb \sr[0]~5 (
	.dataa(altera_internal_jtag1),
	.datab(sr_1),
	.datac(gnd),
	.datad(\DRsize.000~q ),
	.cin(gnd),
	.combout(\sr[0]~5_combout ),
	.cout());
defparam \sr[0]~5 .lut_mask = 16'hAACC;
defparam \sr[0]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Mux37~0 (
	.dataa(irf_reg_0_2),
	.datab(irf_reg_1_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux37~0_combout ),
	.cout());
defparam \Mux37~0 .lut_mask = 16'h7777;
defparam \Mux37~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~10 (
	.dataa(sr_0),
	.datab(virtual_state_cdr),
	.datac(\the_altera_std_synchronizer2|dreg[0]~q ),
	.datad(\Mux37~0_combout ),
	.cin(gnd),
	.combout(\sr~10_combout ),
	.cout());
defparam \sr~10 .lut_mask = 16'hFFB8;
defparam \sr~10 .sum_lutc_input = "datac";

dffeas \DRsize.100 (
	.clk(altera_internal_jtag),
	.d(\Mux37~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.100~q ),
	.prn(vcc));
defparam \DRsize.100 .is_wysiwyg = "true";
defparam \DRsize.100 .power_up = "low";

cyclone10lp_lcell_comb \sr[35]~6 (
	.dataa(sr_36),
	.datab(altera_internal_jtag1),
	.datac(gnd),
	.datad(\DRsize.100~q ),
	.cin(gnd),
	.combout(\sr[35]~6_combout ),
	.cout());
defparam \sr[35]~6 .lut_mask = 16'hAACC;
defparam \sr[35]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~23 (
	.dataa(sr_35),
	.datab(virtual_state_cdr),
	.datac(irf_reg_0_2),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~23_combout ),
	.cout());
defparam \sr~23 .lut_mask = 16'hFFFE;
defparam \sr~23 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~24 (
	.dataa(state_3),
	.datab(splitter_nodes_receive_1_3),
	.datac(\the_altera_std_synchronizer1|dreg[0]~q ),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\sr~24_combout ),
	.cout());
defparam \sr~24 .lut_mask = 16'hFEFF;
defparam \sr~24 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~25 (
	.dataa(\sr~23_combout ),
	.datab(\sr~24_combout ),
	.datac(irf_reg_0_2),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~25_combout ),
	.cout());
defparam \sr~25 .lut_mask = 16'hEFFF;
defparam \sr~25 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr[31]~50 (
	.dataa(irf_reg_0_2),
	.datab(irf_reg_1_2),
	.datac(break_readreg_30),
	.datad(MonDReg_30),
	.cin(gnd),
	.combout(\sr[31]~50_combout ),
	.cout());
defparam \sr[31]~50 .lut_mask = 16'hFFF6;
defparam \sr[31]~50 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr[31]~7 (
	.dataa(sr_31),
	.datab(virtual_state_cdr),
	.datac(irf_reg_0_2),
	.datad(\sr[31]~50_combout ),
	.cin(gnd),
	.combout(\sr[31]~7_combout ),
	.cout());
defparam \sr[31]~7 .lut_mask = 16'hBF8F;
defparam \sr[31]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Mux30~0 (
	.dataa(break_readreg_6),
	.datab(MonDReg_6),
	.datac(irf_reg_1_2),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\Mux30~0_combout ),
	.cout());
defparam \Mux30~0 .lut_mask = 16'hACFF;
defparam \Mux30~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr[7]~8 (
	.dataa(\Mux30~0_combout ),
	.datab(sr_7),
	.datac(gnd),
	.datad(virtual_state_cdr),
	.cin(gnd),
	.combout(\sr[7]~8_combout ),
	.cout());
defparam \sr[7]~8 .lut_mask = 16'hAACC;
defparam \sr[7]~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr[33]~83 (
	.dataa(irf_reg_0_2),
	.datab(irf_reg_1_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sr[33]~83_combout ),
	.cout());
defparam \sr[33]~83 .lut_mask = 16'hEEEE;
defparam \sr[33]~83 .sum_lutc_input = "datac";

dffeas \DRsize.010 (
	.clk(altera_internal_jtag),
	.d(\sr[33]~83_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.010~q ),
	.prn(vcc));
defparam \DRsize.010 .is_wysiwyg = "true";
defparam \DRsize.010 .power_up = "low";

cyclone10lp_lcell_comb \sr[15]~9 (
	.dataa(sr_16),
	.datab(altera_internal_jtag1),
	.datac(gnd),
	.datad(\DRsize.010~q ),
	.cin(gnd),
	.combout(\sr[15]~9_combout ),
	.cout());
defparam \sr[15]~9 .lut_mask = 16'hAACC;
defparam \sr[15]~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~71 (
	.dataa(break_readreg_14),
	.datab(MonDReg_14),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~71_combout ),
	.cout());
defparam \sr~71 .lut_mask = 16'hAACC;
defparam \sr~71 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~72 (
	.dataa(sr_15),
	.datab(virtual_state_cdr),
	.datac(\sr~71_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~72_combout ),
	.cout());
defparam \sr~72 .lut_mask = 16'hB8FF;
defparam \sr~72 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~11 (
	.dataa(break_readreg_0),
	.datab(MonDReg_0),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~11_combout ),
	.cout());
defparam \sr~11 .lut_mask = 16'hAACC;
defparam \sr~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~12 (
	.dataa(sr_2),
	.datab(virtual_state_sdr),
	.datac(\sr~11_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~12_combout ),
	.cout());
defparam \sr~12 .lut_mask = 16'hB8FF;
defparam \sr~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr[13]~13 (
	.dataa(splitter_nodes_receive_1_3),
	.datab(state_3),
	.datac(state_4),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\sr[13]~13_combout ),
	.cout());
defparam \sr[13]~13 .lut_mask = 16'hFEFF;
defparam \sr[13]~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~14 (
	.dataa(break_readreg_1),
	.datab(MonDReg_1),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~14_combout ),
	.cout());
defparam \sr~14 .lut_mask = 16'hAACC;
defparam \sr~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~15 (
	.dataa(sr_3),
	.datab(virtual_state_sdr),
	.datac(\sr~14_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~15_combout ),
	.cout());
defparam \sr~15 .lut_mask = 16'hB8FF;
defparam \sr~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~16 (
	.dataa(break_readreg_2),
	.datab(MonDReg_2),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~16_combout ),
	.cout());
defparam \sr~16 .lut_mask = 16'hAACC;
defparam \sr~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~17 (
	.dataa(sr_4),
	.datab(virtual_state_sdr),
	.datac(\sr~16_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~17_combout ),
	.cout());
defparam \sr~17 .lut_mask = 16'hB8FF;
defparam \sr~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~18 (
	.dataa(break_readreg_3),
	.datab(MonDReg_3),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~18_combout ),
	.cout());
defparam \sr~18 .lut_mask = 16'hAACC;
defparam \sr~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~19 (
	.dataa(sr_5),
	.datab(virtual_state_sdr),
	.datac(\sr~18_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~19_combout ),
	.cout());
defparam \sr~19 .lut_mask = 16'hB8FF;
defparam \sr~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~20 (
	.dataa(splitter_nodes_receive_1_3),
	.datab(state_4),
	.datac(sr_37),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\sr~20_combout ),
	.cout());
defparam \sr~20 .lut_mask = 16'hFEFF;
defparam \sr~20 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr[36]~21 (
	.dataa(virtual_state_cdr),
	.datab(irf_reg_0_2),
	.datac(irf_reg_1_2),
	.datad(virtual_state_sdr),
	.cin(gnd),
	.combout(\sr[36]~21_combout ),
	.cout());
defparam \sr[36]~21 .lut_mask = 16'hFF7D;
defparam \sr[36]~21 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~22 (
	.dataa(altera_internal_jtag1),
	.datab(splitter_nodes_receive_1_3),
	.datac(state_4),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\sr~22_combout ),
	.cout());
defparam \sr~22 .lut_mask = 16'hFEFF;
defparam \sr~22 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~26 (
	.dataa(break_readreg_16),
	.datab(MonDReg_16),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~26_combout ),
	.cout());
defparam \sr~26 .lut_mask = 16'hAACC;
defparam \sr~26 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~27 (
	.dataa(virtual_state_sdr),
	.datab(irf_reg_0_2),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~27_combout ),
	.cout());
defparam \sr~27 .lut_mask = 16'hEEFF;
defparam \sr~27 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~28 (
	.dataa(virtual_state_sdr),
	.datab(sr_18),
	.datac(\sr~26_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~28_combout ),
	.cout());
defparam \sr~28 .lut_mask = 16'hFEFF;
defparam \sr~28 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr[33]~29 (
	.dataa(virtual_state_cdr),
	.datab(irf_reg_0_2),
	.datac(irf_reg_1_2),
	.datad(virtual_state_sdr),
	.cin(gnd),
	.combout(\sr[33]~29_combout ),
	.cout());
defparam \sr[33]~29 .lut_mask = 16'hFF7F;
defparam \sr[33]~29 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~30 (
	.dataa(sr_35),
	.datab(virtual_state_sdr),
	.datac(monitor_error),
	.datad(\Mux37~0_combout ),
	.cin(gnd),
	.combout(\sr~30_combout ),
	.cout());
defparam \sr~30 .lut_mask = 16'hFFB8;
defparam \sr~30 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~31 (
	.dataa(break_readreg_4),
	.datab(MonDReg_4),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~31_combout ),
	.cout());
defparam \sr~31 .lut_mask = 16'hAACC;
defparam \sr~31 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~32 (
	.dataa(sr_6),
	.datab(virtual_state_sdr),
	.datac(\sr~31_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~32_combout ),
	.cout());
defparam \sr~32 .lut_mask = 16'hB8FF;
defparam \sr~32 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~33 (
	.dataa(break_readreg_25),
	.datab(MonDReg_25),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~33_combout ),
	.cout());
defparam \sr~33 .lut_mask = 16'hAACC;
defparam \sr~33 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~34 (
	.dataa(virtual_state_sdr),
	.datab(sr_27),
	.datac(\sr~33_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~34_combout ),
	.cout());
defparam \sr~34 .lut_mask = 16'hFEFF;
defparam \sr~34 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~35 (
	.dataa(break_readreg_27),
	.datab(MonDReg_27),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~35_combout ),
	.cout());
defparam \sr~35 .lut_mask = 16'hAACC;
defparam \sr~35 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~36 (
	.dataa(virtual_state_sdr),
	.datab(sr_29),
	.datac(\sr~35_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~36_combout ),
	.cout());
defparam \sr~36 .lut_mask = 16'hFEFF;
defparam \sr~36 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~37 (
	.dataa(break_readreg_26),
	.datab(MonDReg_26),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~37_combout ),
	.cout());
defparam \sr~37 .lut_mask = 16'hAACC;
defparam \sr~37 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~38 (
	.dataa(virtual_state_sdr),
	.datab(sr_28),
	.datac(\sr~37_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~38_combout ),
	.cout());
defparam \sr~38 .lut_mask = 16'hFEFF;
defparam \sr~38 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~39 (
	.dataa(break_readreg_24),
	.datab(MonDReg_24),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~39_combout ),
	.cout());
defparam \sr~39 .lut_mask = 16'hAACC;
defparam \sr~39 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~40 (
	.dataa(virtual_state_sdr),
	.datab(sr_26),
	.datac(\sr~39_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~40_combout ),
	.cout());
defparam \sr~40 .lut_mask = 16'hFEFF;
defparam \sr~40 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~41 (
	.dataa(break_readreg_20),
	.datab(MonDReg_20),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~41_combout ),
	.cout());
defparam \sr~41 .lut_mask = 16'hAACC;
defparam \sr~41 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~42 (
	.dataa(virtual_state_sdr),
	.datab(sr_22),
	.datac(\sr~41_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~42_combout ),
	.cout());
defparam \sr~42 .lut_mask = 16'hFEFF;
defparam \sr~42 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~43 (
	.dataa(break_readreg_19),
	.datab(MonDReg_19),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~43_combout ),
	.cout());
defparam \sr~43 .lut_mask = 16'hAACC;
defparam \sr~43 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~44 (
	.dataa(virtual_state_sdr),
	.datab(sr_21),
	.datac(\sr~43_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~44_combout ),
	.cout());
defparam \sr~44 .lut_mask = 16'hFEFF;
defparam \sr~44 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~45 (
	.dataa(break_readreg_17),
	.datab(MonDReg_17),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~45_combout ),
	.cout());
defparam \sr~45 .lut_mask = 16'hAACC;
defparam \sr~45 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~46 (
	.dataa(virtual_state_sdr),
	.datab(sr_19),
	.datac(\sr~45_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~46_combout ),
	.cout());
defparam \sr~46 .lut_mask = 16'hFEFF;
defparam \sr~46 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~47 (
	.dataa(sr_34),
	.datab(virtual_state_sdr),
	.datac(resetlatch),
	.datad(\Mux37~0_combout ),
	.cin(gnd),
	.combout(\sr~47_combout ),
	.cout());
defparam \sr~47 .lut_mask = 16'hFFB8;
defparam \sr~47 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~48 (
	.dataa(break_readreg_31),
	.datab(MonDReg_31),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~48_combout ),
	.cout());
defparam \sr~48 .lut_mask = 16'hAACC;
defparam \sr~48 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~49 (
	.dataa(virtual_state_sdr),
	.datab(sr_33),
	.datac(\sr~48_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~49_combout ),
	.cout());
defparam \sr~49 .lut_mask = 16'hFEFF;
defparam \sr~49 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~51 (
	.dataa(break_readreg_29),
	.datab(MonDReg_29),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~51_combout ),
	.cout());
defparam \sr~51 .lut_mask = 16'hAACC;
defparam \sr~51 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~52 (
	.dataa(virtual_state_sdr),
	.datab(sr_31),
	.datac(\sr~51_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~52_combout ),
	.cout());
defparam \sr~52 .lut_mask = 16'hFEFF;
defparam \sr~52 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~53 (
	.dataa(break_readreg_28),
	.datab(MonDReg_28),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~53_combout ),
	.cout());
defparam \sr~53 .lut_mask = 16'hAACC;
defparam \sr~53 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~54 (
	.dataa(virtual_state_sdr),
	.datab(sr_30),
	.datac(\sr~53_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~54_combout ),
	.cout());
defparam \sr~54 .lut_mask = 16'hFEFF;
defparam \sr~54 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~55 (
	.dataa(break_readreg_5),
	.datab(MonDReg_5),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~55_combout ),
	.cout());
defparam \sr~55 .lut_mask = 16'hAACC;
defparam \sr~55 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~56 (
	.dataa(sr_7),
	.datab(virtual_state_sdr),
	.datac(\sr~55_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~56_combout ),
	.cout());
defparam \sr~56 .lut_mask = 16'hB8FF;
defparam \sr~56 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~57 (
	.dataa(break_readreg_18),
	.datab(MonDReg_18),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~57_combout ),
	.cout());
defparam \sr~57 .lut_mask = 16'hAACC;
defparam \sr~57 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~58 (
	.dataa(virtual_state_sdr),
	.datab(sr_20),
	.datac(\sr~57_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~58_combout ),
	.cout());
defparam \sr~58 .lut_mask = 16'hFEFF;
defparam \sr~58 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~59 (
	.dataa(break_readreg_21),
	.datab(MonDReg_21),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~59_combout ),
	.cout());
defparam \sr~59 .lut_mask = 16'hAACC;
defparam \sr~59 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~60 (
	.dataa(virtual_state_sdr),
	.datab(sr_23),
	.datac(\sr~59_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~60_combout ),
	.cout());
defparam \sr~60 .lut_mask = 16'hFEFF;
defparam \sr~60 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~61 (
	.dataa(break_readreg_22),
	.datab(MonDReg_22),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~61_combout ),
	.cout());
defparam \sr~61 .lut_mask = 16'hAACC;
defparam \sr~61 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~62 (
	.dataa(virtual_state_sdr),
	.datab(sr_24),
	.datac(\sr~61_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~62_combout ),
	.cout());
defparam \sr~62 .lut_mask = 16'hFEFF;
defparam \sr~62 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~63 (
	.dataa(break_readreg_15),
	.datab(MonDReg_15),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~63_combout ),
	.cout());
defparam \sr~63 .lut_mask = 16'hAACC;
defparam \sr~63 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~64 (
	.dataa(virtual_state_sdr),
	.datab(sr_17),
	.datac(\sr~63_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~64_combout ),
	.cout());
defparam \sr~64 .lut_mask = 16'hFEFF;
defparam \sr~64 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~65 (
	.dataa(break_readreg_7),
	.datab(MonDReg_7),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~65_combout ),
	.cout());
defparam \sr~65 .lut_mask = 16'hAACC;
defparam \sr~65 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~66 (
	.dataa(sr_9),
	.datab(virtual_state_sdr),
	.datac(\sr~65_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~66_combout ),
	.cout());
defparam \sr~66 .lut_mask = 16'hB8FF;
defparam \sr~66 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~67 (
	.dataa(break_readreg_23),
	.datab(MonDReg_23),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~67_combout ),
	.cout());
defparam \sr~67 .lut_mask = 16'hAACC;
defparam \sr~67 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~68 (
	.dataa(virtual_state_sdr),
	.datab(sr_25),
	.datac(\sr~67_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~68_combout ),
	.cout());
defparam \sr~68 .lut_mask = 16'hFEFF;
defparam \sr~68 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~69 (
	.dataa(break_readreg_13),
	.datab(MonDReg_13),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~69_combout ),
	.cout());
defparam \sr~69 .lut_mask = 16'hAACC;
defparam \sr~69 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~70 (
	.dataa(sr_15),
	.datab(virtual_state_sdr),
	.datac(\sr~69_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~70_combout ),
	.cout());
defparam \sr~70 .lut_mask = 16'hB8FF;
defparam \sr~70 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~73 (
	.dataa(break_readreg_12),
	.datab(MonDReg_12),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~73_combout ),
	.cout());
defparam \sr~73 .lut_mask = 16'hAACC;
defparam \sr~73 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~74 (
	.dataa(sr_14),
	.datab(virtual_state_sdr),
	.datac(\sr~73_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~74_combout ),
	.cout());
defparam \sr~74 .lut_mask = 16'hB8FF;
defparam \sr~74 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~75 (
	.dataa(break_readreg_11),
	.datab(MonDReg_11),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~75_combout ),
	.cout());
defparam \sr~75 .lut_mask = 16'hAACC;
defparam \sr~75 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~76 (
	.dataa(sr_13),
	.datab(virtual_state_sdr),
	.datac(\sr~75_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~76_combout ),
	.cout());
defparam \sr~76 .lut_mask = 16'hB8FF;
defparam \sr~76 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~77 (
	.dataa(break_readreg_10),
	.datab(MonDReg_10),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~77_combout ),
	.cout());
defparam \sr~77 .lut_mask = 16'hAACC;
defparam \sr~77 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~78 (
	.dataa(sr_12),
	.datab(virtual_state_sdr),
	.datac(\sr~77_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~78_combout ),
	.cout());
defparam \sr~78 .lut_mask = 16'hB8FF;
defparam \sr~78 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~79 (
	.dataa(break_readreg_9),
	.datab(MonDReg_9),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~79_combout ),
	.cout());
defparam \sr~79 .lut_mask = 16'hAACC;
defparam \sr~79 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~80 (
	.dataa(sr_11),
	.datab(virtual_state_sdr),
	.datac(\sr~79_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~80_combout ),
	.cout());
defparam \sr~80 .lut_mask = 16'hB8FF;
defparam \sr~80 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~81 (
	.dataa(break_readreg_8),
	.datab(MonDReg_8),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~81_combout ),
	.cout());
defparam \sr~81 .lut_mask = 16'hAACC;
defparam \sr~81 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \sr~82 (
	.dataa(sr_10),
	.datab(virtual_state_sdr),
	.datac(\sr~81_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~82_combout ),
	.cout());
defparam \sr~82 .lut_mask = 16'hB8FF;
defparam \sr~82 .sum_lutc_input = "datac";

endmodule

module processor_altera_std_synchronizer_2 (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module processor_altera_std_synchronizer_3 (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module processor_sld_virtual_jtag_basic_1 (
	virtual_state_cdr1,
	virtual_state_sdr,
	virtual_state_uir,
	virtual_state_udr,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3)/* synthesis synthesis_greybox=1 */;
output 	virtual_state_cdr1;
output 	virtual_state_sdr;
output 	virtual_state_uir;
output 	virtual_state_udr;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclone10lp_lcell_comb virtual_state_cdr(
	.dataa(virtual_ir_scan_reg),
	.datab(gnd),
	.datac(state_3),
	.datad(splitter_nodes_receive_1_3),
	.cin(gnd),
	.combout(virtual_state_cdr1),
	.cout());
defparam virtual_state_cdr.lut_mask = 16'hAFFF;
defparam virtual_state_cdr.sum_lutc_input = "datac";

cyclone10lp_lcell_comb \virtual_state_sdr~0 (
	.dataa(splitter_nodes_receive_1_3),
	.datab(state_4),
	.datac(gnd),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(virtual_state_sdr),
	.cout());
defparam \virtual_state_sdr~0 .lut_mask = 16'hEEFF;
defparam \virtual_state_sdr~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \virtual_state_uir~0 (
	.dataa(virtual_ir_scan_reg),
	.datab(splitter_nodes_receive_1_3),
	.datac(state_8),
	.datad(gnd),
	.cin(gnd),
	.combout(virtual_state_uir),
	.cout());
defparam \virtual_state_uir~0 .lut_mask = 16'hFEFE;
defparam \virtual_state_uir~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \virtual_state_udr~0 (
	.dataa(splitter_nodes_receive_1_3),
	.datab(state_8),
	.datac(gnd),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(virtual_state_udr),
	.cout());
defparam \virtual_state_udr~0 .lut_mask = 16'hEEFF;
defparam \virtual_state_udr~0 .sum_lutc_input = "datac";

endmodule

module processor_processor_nios2_gen2_0_cpu_nios2_avalon_reg (
	r_sync_rst,
	write,
	address_8,
	debugaccess,
	writedata_0,
	address_0,
	address_1,
	address_2,
	address_3,
	address_4,
	address_5,
	address_6,
	address_7,
	Equal0,
	take_action_ocireg,
	oci_ienable_0,
	oci_ienable_1,
	oci_single_step_mode1,
	writedata_1,
	Equal1,
	writedata_3,
	oci_ienable_31,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	write;
input 	address_8;
input 	debugaccess;
input 	writedata_0;
input 	address_0;
input 	address_1;
input 	address_2;
input 	address_3;
input 	address_4;
input 	address_5;
input 	address_6;
input 	address_7;
output 	Equal0;
output 	take_action_ocireg;
output 	oci_ienable_0;
output 	oci_ienable_1;
output 	oci_single_step_mode1;
input 	writedata_1;
output 	Equal1;
input 	writedata_3;
output 	oci_ienable_31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \oci_ienable[0]~0_combout ;
wire \take_action_oci_intr_mask_reg~0_combout ;
wire \oci_ienable[1]~1_combout ;
wire \oci_single_step_mode~0_combout ;


cyclone10lp_lcell_comb \Equal0~2 (
	.dataa(\Equal0~0_combout ),
	.datab(\Equal0~1_combout ),
	.datac(gnd),
	.datad(address_0),
	.cin(gnd),
	.combout(Equal0),
	.cout());
defparam \Equal0~2 .lut_mask = 16'hEEFF;
defparam \Equal0~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \take_action_ocireg~0 (
	.dataa(write),
	.datab(debugaccess),
	.datac(Equal0),
	.datad(gnd),
	.cin(gnd),
	.combout(take_action_ocireg),
	.cout());
defparam \take_action_ocireg~0 .lut_mask = 16'hFEFE;
defparam \take_action_ocireg~0 .sum_lutc_input = "datac";

dffeas \oci_ienable[0] (
	.clk(clk_clk),
	.d(\oci_ienable[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_action_oci_intr_mask_reg~0_combout ),
	.q(oci_ienable_0),
	.prn(vcc));
defparam \oci_ienable[0] .is_wysiwyg = "true";
defparam \oci_ienable[0] .power_up = "low";

dffeas \oci_ienable[1] (
	.clk(clk_clk),
	.d(\oci_ienable[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_action_oci_intr_mask_reg~0_combout ),
	.q(oci_ienable_1),
	.prn(vcc));
defparam \oci_ienable[1] .is_wysiwyg = "true";
defparam \oci_ienable[1] .power_up = "low";

dffeas oci_single_step_mode(
	.clk(clk_clk),
	.d(\oci_single_step_mode~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(oci_single_step_mode1),
	.prn(vcc));
defparam oci_single_step_mode.is_wysiwyg = "true";
defparam oci_single_step_mode.power_up = "low";

cyclone10lp_lcell_comb \Equal1~0 (
	.dataa(address_0),
	.datab(\Equal0~0_combout ),
	.datac(\Equal0~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(Equal1),
	.cout());
defparam \Equal1~0 .lut_mask = 16'hFEFE;
defparam \Equal1~0 .sum_lutc_input = "datac";

dffeas \oci_ienable[31] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_action_oci_intr_mask_reg~0_combout ),
	.q(oci_ienable_31),
	.prn(vcc));
defparam \oci_ienable[31] .is_wysiwyg = "true";
defparam \oci_ienable[31] .power_up = "low";

cyclone10lp_lcell_comb \Equal0~0 (
	.dataa(address_8),
	.datab(address_5),
	.datac(address_6),
	.datad(address_7),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hBFFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal0~1 (
	.dataa(address_1),
	.datab(address_2),
	.datac(address_3),
	.datad(address_4),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'h7FFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \oci_ienable[0]~0 (
	.dataa(writedata_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\oci_ienable[0]~0_combout ),
	.cout());
defparam \oci_ienable[0]~0 .lut_mask = 16'h5555;
defparam \oci_ienable[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \take_action_oci_intr_mask_reg~0 (
	.dataa(write),
	.datab(debugaccess),
	.datac(Equal1),
	.datad(gnd),
	.cin(gnd),
	.combout(\take_action_oci_intr_mask_reg~0_combout ),
	.cout());
defparam \take_action_oci_intr_mask_reg~0 .lut_mask = 16'hFEFE;
defparam \take_action_oci_intr_mask_reg~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \oci_ienable[1]~1 (
	.dataa(writedata_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\oci_ienable[1]~1_combout ),
	.cout());
defparam \oci_ienable[1]~1 .lut_mask = 16'h5555;
defparam \oci_ienable[1]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \oci_single_step_mode~0 (
	.dataa(writedata_3),
	.datab(oci_single_step_mode1),
	.datac(gnd),
	.datad(take_action_ocireg),
	.cin(gnd),
	.combout(\oci_single_step_mode~0_combout ),
	.cout());
defparam \oci_single_step_mode~0 .lut_mask = 16'hAACC;
defparam \oci_single_step_mode~0 .sum_lutc_input = "datac";

endmodule

module processor_processor_nios2_gen2_0_cpu_nios2_oci_break (
	break_readreg_0,
	break_readreg_1,
	jdo_0,
	jdo_36,
	jdo_37,
	ir_0,
	ir_1,
	enable_action_strobe,
	jdo_3,
	jdo_17,
	break_readreg_2,
	jdo_1,
	jdo_4,
	jdo_26,
	jdo_28,
	jdo_27,
	jdo_25,
	jdo_21,
	jdo_20,
	jdo_31,
	jdo_30,
	jdo_29,
	break_readreg_3,
	jdo_2,
	jdo_5,
	jdo_19,
	jdo_18,
	break_readreg_16,
	break_readreg_4,
	jdo_6,
	break_readreg_25,
	break_readreg_27,
	break_readreg_26,
	break_readreg_24,
	break_readreg_20,
	break_readreg_19,
	jdo_23,
	break_readreg_17,
	jdo_16,
	break_readreg_31,
	break_readreg_30,
	break_readreg_29,
	break_readreg_28,
	break_readreg_5,
	jdo_7,
	jdo_24,
	break_readreg_18,
	break_readreg_21,
	jdo_22,
	jdo_8,
	jdo_14,
	jdo_15,
	jdo_13,
	jdo_12,
	jdo_11,
	jdo_10,
	jdo_9,
	break_readreg_6,
	break_readreg_22,
	break_readreg_15,
	break_readreg_7,
	break_readreg_23,
	break_readreg_13,
	break_readreg_14,
	break_readreg_12,
	break_readreg_11,
	break_readreg_10,
	break_readreg_9,
	break_readreg_8,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	break_readreg_0;
output 	break_readreg_1;
input 	jdo_0;
input 	jdo_36;
input 	jdo_37;
input 	ir_0;
input 	ir_1;
input 	enable_action_strobe;
input 	jdo_3;
input 	jdo_17;
output 	break_readreg_2;
input 	jdo_1;
input 	jdo_4;
input 	jdo_26;
input 	jdo_28;
input 	jdo_27;
input 	jdo_25;
input 	jdo_21;
input 	jdo_20;
input 	jdo_31;
input 	jdo_30;
input 	jdo_29;
output 	break_readreg_3;
input 	jdo_2;
input 	jdo_5;
input 	jdo_19;
input 	jdo_18;
output 	break_readreg_16;
output 	break_readreg_4;
input 	jdo_6;
output 	break_readreg_25;
output 	break_readreg_27;
output 	break_readreg_26;
output 	break_readreg_24;
output 	break_readreg_20;
output 	break_readreg_19;
input 	jdo_23;
output 	break_readreg_17;
input 	jdo_16;
output 	break_readreg_31;
output 	break_readreg_30;
output 	break_readreg_29;
output 	break_readreg_28;
output 	break_readreg_5;
input 	jdo_7;
input 	jdo_24;
output 	break_readreg_18;
output 	break_readreg_21;
input 	jdo_22;
input 	jdo_8;
input 	jdo_14;
input 	jdo_15;
input 	jdo_13;
input 	jdo_12;
input 	jdo_11;
input 	jdo_10;
input 	jdo_9;
output 	break_readreg_6;
output 	break_readreg_22;
output 	break_readreg_15;
output 	break_readreg_7;
output 	break_readreg_23;
output 	break_readreg_13;
output 	break_readreg_14;
output 	break_readreg_12;
output 	break_readreg_11;
output 	break_readreg_10;
output 	break_readreg_9;
output 	break_readreg_8;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \break_readreg~0_combout ;
wire \break_readreg[19]~1_combout ;
wire \break_readreg~2_combout ;
wire \break_readreg~3_combout ;
wire \break_readreg~4_combout ;
wire \break_readreg~5_combout ;
wire \break_readreg~6_combout ;
wire \break_readreg~7_combout ;
wire \break_readreg~8_combout ;
wire \break_readreg~9_combout ;
wire \break_readreg~10_combout ;
wire \break_readreg~11_combout ;
wire \break_readreg~12_combout ;
wire \break_readreg~13_combout ;
wire \break_readreg~14_combout ;
wire \break_readreg~15_combout ;
wire \break_readreg~16_combout ;
wire \break_readreg~17_combout ;
wire \break_readreg~18_combout ;
wire \break_readreg~19_combout ;
wire \break_readreg~20_combout ;
wire \break_readreg~21_combout ;
wire \break_readreg~22_combout ;
wire \break_readreg~23_combout ;
wire \break_readreg~24_combout ;
wire \break_readreg~25_combout ;
wire \break_readreg~26_combout ;
wire \break_readreg~27_combout ;
wire \break_readreg~28_combout ;
wire \break_readreg~29_combout ;
wire \break_readreg~30_combout ;
wire \break_readreg~31_combout ;
wire \break_readreg~32_combout ;


dffeas \break_readreg[0] (
	.clk(clk_clk),
	.d(\break_readreg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_0),
	.prn(vcc));
defparam \break_readreg[0] .is_wysiwyg = "true";
defparam \break_readreg[0] .power_up = "low";

dffeas \break_readreg[1] (
	.clk(clk_clk),
	.d(\break_readreg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_1),
	.prn(vcc));
defparam \break_readreg[1] .is_wysiwyg = "true";
defparam \break_readreg[1] .power_up = "low";

dffeas \break_readreg[2] (
	.clk(clk_clk),
	.d(\break_readreg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_2),
	.prn(vcc));
defparam \break_readreg[2] .is_wysiwyg = "true";
defparam \break_readreg[2] .power_up = "low";

dffeas \break_readreg[3] (
	.clk(clk_clk),
	.d(\break_readreg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_3),
	.prn(vcc));
defparam \break_readreg[3] .is_wysiwyg = "true";
defparam \break_readreg[3] .power_up = "low";

dffeas \break_readreg[16] (
	.clk(clk_clk),
	.d(\break_readreg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_16),
	.prn(vcc));
defparam \break_readreg[16] .is_wysiwyg = "true";
defparam \break_readreg[16] .power_up = "low";

dffeas \break_readreg[4] (
	.clk(clk_clk),
	.d(\break_readreg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_4),
	.prn(vcc));
defparam \break_readreg[4] .is_wysiwyg = "true";
defparam \break_readreg[4] .power_up = "low";

dffeas \break_readreg[25] (
	.clk(clk_clk),
	.d(\break_readreg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_25),
	.prn(vcc));
defparam \break_readreg[25] .is_wysiwyg = "true";
defparam \break_readreg[25] .power_up = "low";

dffeas \break_readreg[27] (
	.clk(clk_clk),
	.d(\break_readreg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_27),
	.prn(vcc));
defparam \break_readreg[27] .is_wysiwyg = "true";
defparam \break_readreg[27] .power_up = "low";

dffeas \break_readreg[26] (
	.clk(clk_clk),
	.d(\break_readreg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_26),
	.prn(vcc));
defparam \break_readreg[26] .is_wysiwyg = "true";
defparam \break_readreg[26] .power_up = "low";

dffeas \break_readreg[24] (
	.clk(clk_clk),
	.d(\break_readreg~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_24),
	.prn(vcc));
defparam \break_readreg[24] .is_wysiwyg = "true";
defparam \break_readreg[24] .power_up = "low";

dffeas \break_readreg[20] (
	.clk(clk_clk),
	.d(\break_readreg~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_20),
	.prn(vcc));
defparam \break_readreg[20] .is_wysiwyg = "true";
defparam \break_readreg[20] .power_up = "low";

dffeas \break_readreg[19] (
	.clk(clk_clk),
	.d(\break_readreg~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_19),
	.prn(vcc));
defparam \break_readreg[19] .is_wysiwyg = "true";
defparam \break_readreg[19] .power_up = "low";

dffeas \break_readreg[17] (
	.clk(clk_clk),
	.d(\break_readreg~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_17),
	.prn(vcc));
defparam \break_readreg[17] .is_wysiwyg = "true";
defparam \break_readreg[17] .power_up = "low";

dffeas \break_readreg[31] (
	.clk(clk_clk),
	.d(\break_readreg~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_31),
	.prn(vcc));
defparam \break_readreg[31] .is_wysiwyg = "true";
defparam \break_readreg[31] .power_up = "low";

dffeas \break_readreg[30] (
	.clk(clk_clk),
	.d(\break_readreg~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_30),
	.prn(vcc));
defparam \break_readreg[30] .is_wysiwyg = "true";
defparam \break_readreg[30] .power_up = "low";

dffeas \break_readreg[29] (
	.clk(clk_clk),
	.d(\break_readreg~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_29),
	.prn(vcc));
defparam \break_readreg[29] .is_wysiwyg = "true";
defparam \break_readreg[29] .power_up = "low";

dffeas \break_readreg[28] (
	.clk(clk_clk),
	.d(\break_readreg~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_28),
	.prn(vcc));
defparam \break_readreg[28] .is_wysiwyg = "true";
defparam \break_readreg[28] .power_up = "low";

dffeas \break_readreg[5] (
	.clk(clk_clk),
	.d(\break_readreg~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_5),
	.prn(vcc));
defparam \break_readreg[5] .is_wysiwyg = "true";
defparam \break_readreg[5] .power_up = "low";

dffeas \break_readreg[18] (
	.clk(clk_clk),
	.d(\break_readreg~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_18),
	.prn(vcc));
defparam \break_readreg[18] .is_wysiwyg = "true";
defparam \break_readreg[18] .power_up = "low";

dffeas \break_readreg[21] (
	.clk(clk_clk),
	.d(\break_readreg~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_21),
	.prn(vcc));
defparam \break_readreg[21] .is_wysiwyg = "true";
defparam \break_readreg[21] .power_up = "low";

dffeas \break_readreg[6] (
	.clk(clk_clk),
	.d(\break_readreg~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_6),
	.prn(vcc));
defparam \break_readreg[6] .is_wysiwyg = "true";
defparam \break_readreg[6] .power_up = "low";

dffeas \break_readreg[22] (
	.clk(clk_clk),
	.d(\break_readreg~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_22),
	.prn(vcc));
defparam \break_readreg[22] .is_wysiwyg = "true";
defparam \break_readreg[22] .power_up = "low";

dffeas \break_readreg[15] (
	.clk(clk_clk),
	.d(\break_readreg~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_15),
	.prn(vcc));
defparam \break_readreg[15] .is_wysiwyg = "true";
defparam \break_readreg[15] .power_up = "low";

dffeas \break_readreg[7] (
	.clk(clk_clk),
	.d(\break_readreg~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_7),
	.prn(vcc));
defparam \break_readreg[7] .is_wysiwyg = "true";
defparam \break_readreg[7] .power_up = "low";

dffeas \break_readreg[23] (
	.clk(clk_clk),
	.d(\break_readreg~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_23),
	.prn(vcc));
defparam \break_readreg[23] .is_wysiwyg = "true";
defparam \break_readreg[23] .power_up = "low";

dffeas \break_readreg[13] (
	.clk(clk_clk),
	.d(\break_readreg~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_13),
	.prn(vcc));
defparam \break_readreg[13] .is_wysiwyg = "true";
defparam \break_readreg[13] .power_up = "low";

dffeas \break_readreg[14] (
	.clk(clk_clk),
	.d(\break_readreg~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_14),
	.prn(vcc));
defparam \break_readreg[14] .is_wysiwyg = "true";
defparam \break_readreg[14] .power_up = "low";

dffeas \break_readreg[12] (
	.clk(clk_clk),
	.d(\break_readreg~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_12),
	.prn(vcc));
defparam \break_readreg[12] .is_wysiwyg = "true";
defparam \break_readreg[12] .power_up = "low";

dffeas \break_readreg[11] (
	.clk(clk_clk),
	.d(\break_readreg~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_11),
	.prn(vcc));
defparam \break_readreg[11] .is_wysiwyg = "true";
defparam \break_readreg[11] .power_up = "low";

dffeas \break_readreg[10] (
	.clk(clk_clk),
	.d(\break_readreg~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_10),
	.prn(vcc));
defparam \break_readreg[10] .is_wysiwyg = "true";
defparam \break_readreg[10] .power_up = "low";

dffeas \break_readreg[9] (
	.clk(clk_clk),
	.d(\break_readreg~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_9),
	.prn(vcc));
defparam \break_readreg[9] .is_wysiwyg = "true";
defparam \break_readreg[9] .power_up = "low";

dffeas \break_readreg[8] (
	.clk(clk_clk),
	.d(\break_readreg~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_8),
	.prn(vcc));
defparam \break_readreg[8] .is_wysiwyg = "true";
defparam \break_readreg[8] .power_up = "low";

cyclone10lp_lcell_comb \break_readreg~0 (
	.dataa(jdo_0),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(gnd),
	.cin(gnd),
	.combout(\break_readreg~0_combout ),
	.cout());
defparam \break_readreg~0 .lut_mask = 16'hFEFE;
defparam \break_readreg~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg[19]~1 (
	.dataa(ir_0),
	.datab(gnd),
	.datac(ir_1),
	.datad(enable_action_strobe),
	.cin(gnd),
	.combout(\break_readreg[19]~1_combout ),
	.cout());
defparam \break_readreg[19]~1 .lut_mask = 16'hFFF5;
defparam \break_readreg[19]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg~2 (
	.dataa(jdo_1),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(gnd),
	.cin(gnd),
	.combout(\break_readreg~2_combout ),
	.cout());
defparam \break_readreg~2 .lut_mask = 16'hFEFE;
defparam \break_readreg~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg~3 (
	.dataa(jdo_2),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(gnd),
	.cin(gnd),
	.combout(\break_readreg~3_combout ),
	.cout());
defparam \break_readreg~3 .lut_mask = 16'hFEFE;
defparam \break_readreg~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg~4 (
	.dataa(jdo_3),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~4_combout ),
	.cout());
defparam \break_readreg~4 .lut_mask = 16'hFEFF;
defparam \break_readreg~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg~5 (
	.dataa(jdo_16),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~5_combout ),
	.cout());
defparam \break_readreg~5 .lut_mask = 16'hFEFF;
defparam \break_readreg~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg~6 (
	.dataa(jdo_4),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~6_combout ),
	.cout());
defparam \break_readreg~6 .lut_mask = 16'hFEFF;
defparam \break_readreg~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg~7 (
	.dataa(jdo_25),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~7_combout ),
	.cout());
defparam \break_readreg~7 .lut_mask = 16'hFEFF;
defparam \break_readreg~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg~8 (
	.dataa(jdo_27),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~8_combout ),
	.cout());
defparam \break_readreg~8 .lut_mask = 16'hFEFF;
defparam \break_readreg~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg~9 (
	.dataa(jdo_26),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~9_combout ),
	.cout());
defparam \break_readreg~9 .lut_mask = 16'hFEFF;
defparam \break_readreg~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg~10 (
	.dataa(jdo_24),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~10_combout ),
	.cout());
defparam \break_readreg~10 .lut_mask = 16'hFEFF;
defparam \break_readreg~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg~11 (
	.dataa(jdo_20),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~11_combout ),
	.cout());
defparam \break_readreg~11 .lut_mask = 16'hFEFF;
defparam \break_readreg~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg~12 (
	.dataa(jdo_19),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~12_combout ),
	.cout());
defparam \break_readreg~12 .lut_mask = 16'hFEFF;
defparam \break_readreg~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg~13 (
	.dataa(jdo_17),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~13_combout ),
	.cout());
defparam \break_readreg~13 .lut_mask = 16'hFEFF;
defparam \break_readreg~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg~14 (
	.dataa(jdo_31),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~14_combout ),
	.cout());
defparam \break_readreg~14 .lut_mask = 16'hFEFF;
defparam \break_readreg~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg~15 (
	.dataa(jdo_30),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~15_combout ),
	.cout());
defparam \break_readreg~15 .lut_mask = 16'hFEFF;
defparam \break_readreg~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg~16 (
	.dataa(jdo_29),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~16_combout ),
	.cout());
defparam \break_readreg~16 .lut_mask = 16'hFEFF;
defparam \break_readreg~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg~17 (
	.dataa(jdo_28),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~17_combout ),
	.cout());
defparam \break_readreg~17 .lut_mask = 16'hFEFF;
defparam \break_readreg~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg~18 (
	.dataa(jdo_5),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~18_combout ),
	.cout());
defparam \break_readreg~18 .lut_mask = 16'hFEFF;
defparam \break_readreg~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg~19 (
	.dataa(jdo_18),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~19_combout ),
	.cout());
defparam \break_readreg~19 .lut_mask = 16'hFEFF;
defparam \break_readreg~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg~20 (
	.dataa(jdo_21),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~20_combout ),
	.cout());
defparam \break_readreg~20 .lut_mask = 16'hFEFF;
defparam \break_readreg~20 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg~21 (
	.dataa(jdo_6),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~21_combout ),
	.cout());
defparam \break_readreg~21 .lut_mask = 16'hFEFF;
defparam \break_readreg~21 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg~22 (
	.dataa(jdo_22),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~22_combout ),
	.cout());
defparam \break_readreg~22 .lut_mask = 16'hFEFF;
defparam \break_readreg~22 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg~23 (
	.dataa(jdo_15),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~23_combout ),
	.cout());
defparam \break_readreg~23 .lut_mask = 16'hFEFF;
defparam \break_readreg~23 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg~24 (
	.dataa(jdo_7),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~24_combout ),
	.cout());
defparam \break_readreg~24 .lut_mask = 16'hFEFF;
defparam \break_readreg~24 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg~25 (
	.dataa(jdo_23),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~25_combout ),
	.cout());
defparam \break_readreg~25 .lut_mask = 16'hFEFF;
defparam \break_readreg~25 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg~26 (
	.dataa(jdo_13),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~26_combout ),
	.cout());
defparam \break_readreg~26 .lut_mask = 16'hFEFF;
defparam \break_readreg~26 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg~27 (
	.dataa(jdo_14),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~27_combout ),
	.cout());
defparam \break_readreg~27 .lut_mask = 16'hFEFF;
defparam \break_readreg~27 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg~28 (
	.dataa(jdo_12),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~28_combout ),
	.cout());
defparam \break_readreg~28 .lut_mask = 16'hFEFF;
defparam \break_readreg~28 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg~29 (
	.dataa(jdo_11),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~29_combout ),
	.cout());
defparam \break_readreg~29 .lut_mask = 16'hFEFF;
defparam \break_readreg~29 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg~30 (
	.dataa(jdo_10),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~30_combout ),
	.cout());
defparam \break_readreg~30 .lut_mask = 16'hFEFF;
defparam \break_readreg~30 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg~31 (
	.dataa(jdo_9),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~31_combout ),
	.cout());
defparam \break_readreg~31 .lut_mask = 16'hFEFF;
defparam \break_readreg~31 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_readreg~32 (
	.dataa(jdo_8),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~32_combout ),
	.cout());
defparam \break_readreg~32 .lut_mask = 16'hFEFF;
defparam \break_readreg~32 .sum_lutc_input = "datac";

endmodule

module processor_processor_nios2_gen2_0_cpu_nios2_oci_debug (
	jtag_break1,
	r_sync_rst,
	monitor_ready1,
	take_action_ocimem_a,
	jdo_34,
	writedata_0,
	take_action_ocireg,
	jdo_25,
	jdo_21,
	jdo_20,
	take_action_ocimem_a1,
	writedata_1,
	monitor_error1,
	jdo_19,
	jdo_18,
	monitor_go1,
	jdo_23,
	resetlatch1,
	jdo_24,
	state_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	jtag_break1;
input 	r_sync_rst;
output 	monitor_ready1;
input 	take_action_ocimem_a;
input 	jdo_34;
input 	writedata_0;
input 	take_action_ocireg;
input 	jdo_25;
input 	jdo_21;
input 	jdo_20;
input 	take_action_ocimem_a1;
input 	writedata_1;
output 	monitor_error1;
input 	jdo_19;
input 	jdo_18;
output 	monitor_go1;
input 	jdo_23;
output 	resetlatch1;
input 	jdo_24;
input 	state_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer|dreg[0]~q ;
wire \break_on_reset~0_combout ;
wire \break_on_reset~q ;
wire \jtag_break~0_combout ;
wire \jtag_break~1_combout ;
wire \always1~0_combout ;
wire \monitor_ready~0_combout ;
wire \monitor_error~0_combout ;
wire \monitor_go~0_combout ;
wire \resetlatch~0_combout ;


processor_altera_std_synchronizer_4 the_altera_std_synchronizer(
	.din(r_sync_rst),
	.dreg_0(\the_altera_std_synchronizer|dreg[0]~q ),
	.clk(clk_clk));

dffeas jtag_break(
	.clk(clk_clk),
	.d(\jtag_break~0_combout ),
	.asdata(\jtag_break~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(vcc),
	.q(jtag_break1),
	.prn(vcc));
defparam jtag_break.is_wysiwyg = "true";
defparam jtag_break.power_up = "low";

dffeas monitor_ready(
	.clk(clk_clk),
	.d(\monitor_ready~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_ready1),
	.prn(vcc));
defparam monitor_ready.is_wysiwyg = "true";
defparam monitor_ready.power_up = "low";

dffeas monitor_error(
	.clk(clk_clk),
	.d(\monitor_error~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_error1),
	.prn(vcc));
defparam monitor_error.is_wysiwyg = "true";
defparam monitor_error.power_up = "low";

dffeas monitor_go(
	.clk(clk_clk),
	.d(\monitor_go~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_go1),
	.prn(vcc));
defparam monitor_go.is_wysiwyg = "true";
defparam monitor_go.power_up = "low";

dffeas resetlatch(
	.clk(clk_clk),
	.d(\resetlatch~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(resetlatch1),
	.prn(vcc));
defparam resetlatch.is_wysiwyg = "true";
defparam resetlatch.power_up = "low";

cyclone10lp_lcell_comb \break_on_reset~0 (
	.dataa(jdo_19),
	.datab(\break_on_reset~q ),
	.datac(take_action_ocimem_a1),
	.datad(jdo_18),
	.cin(gnd),
	.combout(\break_on_reset~0_combout ),
	.cout());
defparam \break_on_reset~0 .lut_mask = 16'hACFF;
defparam \break_on_reset~0 .sum_lutc_input = "datac";

dffeas break_on_reset(
	.clk(clk_clk),
	.d(\break_on_reset~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\break_on_reset~q ),
	.prn(vcc));
defparam break_on_reset.is_wysiwyg = "true";
defparam break_on_reset.power_up = "low";

cyclone10lp_lcell_comb \jtag_break~0 (
	.dataa(jtag_break1),
	.datab(\break_on_reset~q ),
	.datac(gnd),
	.datad(\the_altera_std_synchronizer|dreg[0]~q ),
	.cin(gnd),
	.combout(\jtag_break~0_combout ),
	.cout());
defparam \jtag_break~0 .lut_mask = 16'hAACC;
defparam \jtag_break~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \jtag_break~1 (
	.dataa(jdo_21),
	.datab(jtag_break1),
	.datac(gnd),
	.datad(jdo_20),
	.cin(gnd),
	.combout(\jtag_break~1_combout ),
	.cout());
defparam \jtag_break~1 .lut_mask = 16'hEEFF;
defparam \jtag_break~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \always1~0 (
	.dataa(take_action_ocimem_a),
	.datab(jdo_34),
	.datac(jdo_25),
	.datad(gnd),
	.cin(gnd),
	.combout(\always1~0_combout ),
	.cout());
defparam \always1~0 .lut_mask = 16'hFEFE;
defparam \always1~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \monitor_ready~0 (
	.dataa(monitor_ready1),
	.datab(writedata_0),
	.datac(take_action_ocireg),
	.datad(\always1~0_combout ),
	.cin(gnd),
	.combout(\monitor_ready~0_combout ),
	.cout());
defparam \monitor_ready~0 .lut_mask = 16'hFEFF;
defparam \monitor_ready~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \monitor_error~0 (
	.dataa(monitor_error1),
	.datab(take_action_ocireg),
	.datac(writedata_1),
	.datad(\always1~0_combout ),
	.cin(gnd),
	.combout(\monitor_error~0_combout ),
	.cout());
defparam \monitor_error~0 .lut_mask = 16'hFEFF;
defparam \monitor_error~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \monitor_go~0 (
	.dataa(take_action_ocimem_a1),
	.datab(jdo_23),
	.datac(monitor_go1),
	.datad(state_1),
	.cin(gnd),
	.combout(\monitor_go~0_combout ),
	.cout());
defparam \monitor_go~0 .lut_mask = 16'hFEFF;
defparam \monitor_go~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \resetlatch~0 (
	.dataa(resetlatch1),
	.datab(\the_altera_std_synchronizer|dreg[0]~q ),
	.datac(jdo_24),
	.datad(take_action_ocimem_a1),
	.cin(gnd),
	.combout(\resetlatch~0_combout ),
	.cout());
defparam \resetlatch~0 .lut_mask = 16'hEFFF;
defparam \resetlatch~0 .sum_lutc_input = "datac";

endmodule

module processor_altera_std_synchronizer_4 (
	din,
	dreg_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	din;
output 	dreg_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module processor_processor_nios2_gen2_0_cpu_nios2_ocimem (
	MonDReg_0,
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_22,
	q_a_23,
	q_a_24,
	q_a_25,
	q_a_26,
	q_a_4,
	q_a_3,
	q_a_5,
	q_a_14,
	q_a_15,
	q_a_11,
	q_a_13,
	q_a_16,
	q_a_12,
	q_a_10,
	q_a_9,
	q_a_8,
	q_a_7,
	q_a_6,
	q_a_21,
	q_a_20,
	q_a_19,
	q_a_18,
	q_a_17,
	MonDReg_4,
	MonDReg_29,
	MonDReg_5,
	MonDReg_15,
	MonDReg_12,
	q_a_27,
	q_a_28,
	q_a_29,
	q_a_30,
	q_a_31,
	MonDReg_8,
	MonDReg_18,
	waitrequest1,
	write,
	address_8,
	read,
	MonDReg_1,
	jdo_3,
	jdo_35,
	take_action_ocimem_b,
	take_action_ocimem_a,
	jdo_17,
	take_action_ocimem_a1,
	jdo_34,
	MonDReg_2,
	jdo_4,
	jdo_26,
	jdo_28,
	jdo_27,
	debugaccess,
	r_early_rst,
	writedata_0,
	address_0,
	address_1,
	address_2,
	address_3,
	address_4,
	address_5,
	address_6,
	address_7,
	byteenable_0,
	jdo_25,
	jdo_21,
	jdo_20,
	jdo_33,
	jdo_32,
	jdo_31,
	jdo_30,
	jdo_29,
	MonDReg_3,
	jdo_5,
	writedata_1,
	jdo_19,
	jdo_18,
	writedata_3,
	MonDReg_16,
	jdo_6,
	writedata_2,
	MonDReg_25,
	MonDReg_27,
	MonDReg_26,
	MonDReg_24,
	MonDReg_20,
	MonDReg_19,
	MonDReg_22,
	writedata_22,
	byteenable_2,
	MonDReg_23,
	writedata_23,
	writedata_24,
	byteenable_3,
	writedata_25,
	writedata_26,
	writedata_4,
	jdo_23,
	MonDReg_17,
	jdo_16,
	MonDReg_31,
	MonDReg_30,
	MonDReg_28,
	writedata_5,
	MonDReg_14,
	writedata_14,
	byteenable_1,
	writedata_15,
	MonDReg_11,
	writedata_11,
	MonDReg_13,
	writedata_13,
	writedata_16,
	writedata_12,
	MonDReg_10,
	writedata_10,
	MonDReg_9,
	writedata_9,
	writedata_8,
	MonDReg_7,
	writedata_7,
	MonDReg_6,
	writedata_6,
	MonDReg_21,
	writedata_21,
	writedata_20,
	writedata_19,
	writedata_18,
	writedata_17,
	jdo_7,
	jdo_24,
	jdo_22,
	jdo_8,
	jdo_14,
	jdo_15,
	writedata_27,
	writedata_28,
	writedata_29,
	writedata_30,
	writedata_31,
	jdo_13,
	jdo_12,
	jdo_11,
	jdo_10,
	jdo_9,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	MonDReg_0;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_22;
output 	q_a_23;
output 	q_a_24;
output 	q_a_25;
output 	q_a_26;
output 	q_a_4;
output 	q_a_3;
output 	q_a_5;
output 	q_a_14;
output 	q_a_15;
output 	q_a_11;
output 	q_a_13;
output 	q_a_16;
output 	q_a_12;
output 	q_a_10;
output 	q_a_9;
output 	q_a_8;
output 	q_a_7;
output 	q_a_6;
output 	q_a_21;
output 	q_a_20;
output 	q_a_19;
output 	q_a_18;
output 	q_a_17;
output 	MonDReg_4;
output 	MonDReg_29;
output 	MonDReg_5;
output 	MonDReg_15;
output 	MonDReg_12;
output 	q_a_27;
output 	q_a_28;
output 	q_a_29;
output 	q_a_30;
output 	q_a_31;
output 	MonDReg_8;
output 	MonDReg_18;
output 	waitrequest1;
input 	write;
input 	address_8;
input 	read;
output 	MonDReg_1;
input 	jdo_3;
input 	jdo_35;
input 	take_action_ocimem_b;
input 	take_action_ocimem_a;
input 	jdo_17;
input 	take_action_ocimem_a1;
input 	jdo_34;
output 	MonDReg_2;
input 	jdo_4;
input 	jdo_26;
input 	jdo_28;
input 	jdo_27;
input 	debugaccess;
input 	r_early_rst;
input 	writedata_0;
input 	address_0;
input 	address_1;
input 	address_2;
input 	address_3;
input 	address_4;
input 	address_5;
input 	address_6;
input 	address_7;
input 	byteenable_0;
input 	jdo_25;
input 	jdo_21;
input 	jdo_20;
input 	jdo_33;
input 	jdo_32;
input 	jdo_31;
input 	jdo_30;
input 	jdo_29;
output 	MonDReg_3;
input 	jdo_5;
input 	writedata_1;
input 	jdo_19;
input 	jdo_18;
input 	writedata_3;
output 	MonDReg_16;
input 	jdo_6;
input 	writedata_2;
output 	MonDReg_25;
output 	MonDReg_27;
output 	MonDReg_26;
output 	MonDReg_24;
output 	MonDReg_20;
output 	MonDReg_19;
output 	MonDReg_22;
input 	writedata_22;
input 	byteenable_2;
output 	MonDReg_23;
input 	writedata_23;
input 	writedata_24;
input 	byteenable_3;
input 	writedata_25;
input 	writedata_26;
input 	writedata_4;
input 	jdo_23;
output 	MonDReg_17;
input 	jdo_16;
output 	MonDReg_31;
output 	MonDReg_30;
output 	MonDReg_28;
input 	writedata_5;
output 	MonDReg_14;
input 	writedata_14;
input 	byteenable_1;
input 	writedata_15;
output 	MonDReg_11;
input 	writedata_11;
output 	MonDReg_13;
input 	writedata_13;
input 	writedata_16;
input 	writedata_12;
output 	MonDReg_10;
input 	writedata_10;
output 	MonDReg_9;
input 	writedata_9;
input 	writedata_8;
output 	MonDReg_7;
input 	writedata_7;
output 	MonDReg_6;
input 	writedata_6;
output 	MonDReg_21;
input 	writedata_21;
input 	writedata_20;
input 	writedata_19;
input 	writedata_18;
input 	writedata_17;
input 	jdo_7;
input 	jdo_24;
input 	jdo_22;
input 	jdo_8;
input 	jdo_14;
input 	jdo_15;
input 	writedata_27;
input 	writedata_28;
input 	writedata_29;
input 	writedata_30;
input 	writedata_31;
input 	jdo_13;
input 	jdo_12;
input 	jdo_11;
input 	jdo_10;
input 	jdo_9;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ociram_wr_en~0_combout ;
wire \jtag_ram_wr~q ;
wire \ociram_wr_en~1_combout ;
wire \ociram_reset_req~combout ;
wire \ociram_wr_data[0]~0_combout ;
wire \ociram_addr[0]~0_combout ;
wire \ociram_addr[1]~1_combout ;
wire \ociram_addr[2]~2_combout ;
wire \ociram_addr[3]~3_combout ;
wire \ociram_addr[4]~4_combout ;
wire \ociram_addr[5]~5_combout ;
wire \ociram_addr[6]~6_combout ;
wire \ociram_addr[7]~7_combout ;
wire \ociram_byteenable[0]~0_combout ;
wire \ociram_wr_data[1]~1_combout ;
wire \jtag_ram_wr~0_combout ;
wire \ociram_wr_data[2]~2_combout ;
wire \ociram_wr_data[22]~3_combout ;
wire \ociram_byteenable[2]~1_combout ;
wire \ociram_wr_data[23]~4_combout ;
wire \ociram_wr_data[24]~5_combout ;
wire \ociram_byteenable[3]~2_combout ;
wire \ociram_wr_data[25]~6_combout ;
wire \ociram_wr_data[26]~7_combout ;
wire \ociram_wr_data[4]~8_combout ;
wire \ociram_wr_data[3]~9_combout ;
wire \ociram_wr_data[5]~10_combout ;
wire \ociram_wr_data[14]~11_combout ;
wire \ociram_byteenable[1]~3_combout ;
wire \ociram_wr_data[15]~12_combout ;
wire \ociram_wr_data[11]~13_combout ;
wire \ociram_wr_data[13]~14_combout ;
wire \ociram_wr_data[16]~15_combout ;
wire \ociram_wr_data[12]~16_combout ;
wire \ociram_wr_data[10]~17_combout ;
wire \ociram_wr_data[9]~18_combout ;
wire \ociram_wr_data[8]~19_combout ;
wire \ociram_wr_data[7]~20_combout ;
wire \ociram_wr_data[6]~21_combout ;
wire \ociram_wr_data[21]~22_combout ;
wire \ociram_wr_data[20]~23_combout ;
wire \ociram_wr_data[19]~24_combout ;
wire \ociram_wr_data[18]~25_combout ;
wire \ociram_wr_data[17]~26_combout ;
wire \ociram_wr_data[27]~27_combout ;
wire \ociram_wr_data[28]~28_combout ;
wire \ociram_wr_data[29]~29_combout ;
wire \ociram_wr_data[30]~30_combout ;
wire \ociram_wr_data[31]~31_combout ;
wire \MonARegAddrInc[0]~0_combout ;
wire \MonAReg~0_combout ;
wire \MonAReg[2]~q ;
wire \MonARegAddrInc[0]~1 ;
wire \MonARegAddrInc[1]~2_combout ;
wire \MonAReg~2_combout ;
wire \MonAReg[3]~q ;
wire \MonARegAddrInc[1]~3 ;
wire \MonARegAddrInc[2]~4_combout ;
wire \MonAReg~1_combout ;
wire \MonAReg[4]~q ;
wire \Equal0~0_combout ;
wire \jtag_ram_access~0_combout ;
wire \MonAReg[10]~q ;
wire \MonARegAddrInc[2]~5 ;
wire \MonARegAddrInc[3]~6_combout ;
wire \MonAReg~7_combout ;
wire \MonAReg[5]~q ;
wire \MonARegAddrInc[3]~7 ;
wire \MonARegAddrInc[4]~8_combout ;
wire \MonAReg~6_combout ;
wire \MonAReg[6]~q ;
wire \MonARegAddrInc[4]~9 ;
wire \MonARegAddrInc[5]~10_combout ;
wire \MonAReg~5_combout ;
wire \MonAReg[7]~q ;
wire \MonARegAddrInc[5]~11 ;
wire \MonARegAddrInc[6]~12_combout ;
wire \MonAReg~4_combout ;
wire \MonAReg[8]~q ;
wire \MonARegAddrInc[6]~13 ;
wire \MonARegAddrInc[7]~14_combout ;
wire \MonAReg~3_combout ;
wire \MonAReg[9]~q ;
wire \MonARegAddrInc[7]~15 ;
wire \MonARegAddrInc[8]~16_combout ;
wire \jtag_ram_rd~0_combout ;
wire \jtag_ram_rd~1_combout ;
wire \jtag_ram_rd~q ;
wire \jtag_ram_rd_d1~q ;
wire \MonDReg[0]~0_combout ;
wire \jtag_rd~0_combout ;
wire \jtag_rd~q ;
wire \jtag_rd_d1~q ;
wire \MonDReg[0]~8_combout ;
wire \MonDReg[4]~1_combout ;
wire \Equal0~1_combout ;
wire \MonDReg[29]~7_combout ;
wire \Equal0~2_combout ;
wire \MonDReg[5]~2_combout ;
wire \cfgrom_readdata[15]~0_combout ;
wire \MonDReg[15]~3_combout ;
wire \MonDReg[15]~26_combout ;
wire \MonDReg[12]~4_combout ;
wire \cfgrom_readdata[8]~1_combout ;
wire \MonDReg[8]~6_combout ;
wire \Equal0~3_combout ;
wire \MonDReg[18]~5_combout ;
wire \jtag_ram_access~1_combout ;
wire \jtag_ram_access~q ;
wire \waitrequest~0_combout ;
wire \avalon_ociram_readdata_ready~0_combout ;
wire \avalon_ociram_readdata_ready~1_combout ;
wire \avalon_ociram_readdata_ready~q ;
wire \waitrequest~1_combout ;
wire \MonDReg~9_combout ;
wire \MonDReg~10_combout ;
wire \MonDReg~11_combout ;
wire \MonDReg~12_combout ;
wire \MonDReg~13_combout ;
wire \MonDReg~14_combout ;
wire \MonDReg~15_combout ;
wire \MonDReg~16_combout ;
wire \MonDReg~17_combout ;
wire \MonDReg~18_combout ;
wire \MonDReg~19_combout ;
wire \MonDReg~20_combout ;
wire \MonDReg~21_combout ;
wire \MonDReg~22_combout ;
wire \MonDReg~23_combout ;
wire \MonDReg~24_combout ;
wire \MonDReg~25_combout ;
wire \MonDReg~27_combout ;
wire \MonDReg~28_combout ;
wire \MonDReg~29_combout ;
wire \MonDReg~30_combout ;
wire \MonDReg~31_combout ;
wire \MonDReg~32_combout ;
wire \MonDReg~33_combout ;


processor_processor_nios2_gen2_0_cpu_ociram_sp_ram_module processor_nios2_gen2_0_cpu_ociram_sp_ram(
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_22(q_a_22),
	.q_a_23(q_a_23),
	.q_a_24(q_a_24),
	.q_a_25(q_a_25),
	.q_a_26(q_a_26),
	.q_a_4(q_a_4),
	.q_a_3(q_a_3),
	.q_a_5(q_a_5),
	.q_a_14(q_a_14),
	.q_a_15(q_a_15),
	.q_a_11(q_a_11),
	.q_a_13(q_a_13),
	.q_a_16(q_a_16),
	.q_a_12(q_a_12),
	.q_a_10(q_a_10),
	.q_a_9(q_a_9),
	.q_a_8(q_a_8),
	.q_a_7(q_a_7),
	.q_a_6(q_a_6),
	.q_a_21(q_a_21),
	.q_a_20(q_a_20),
	.q_a_19(q_a_19),
	.q_a_18(q_a_18),
	.q_a_17(q_a_17),
	.q_a_27(q_a_27),
	.q_a_28(q_a_28),
	.q_a_29(q_a_29),
	.q_a_30(q_a_30),
	.q_a_31(q_a_31),
	.ociram_wr_en(\ociram_wr_en~1_combout ),
	.ociram_reset_req(\ociram_reset_req~combout ),
	.ociram_wr_data_0(\ociram_wr_data[0]~0_combout ),
	.ociram_addr_0(\ociram_addr[0]~0_combout ),
	.ociram_addr_1(\ociram_addr[1]~1_combout ),
	.ociram_addr_2(\ociram_addr[2]~2_combout ),
	.ociram_addr_3(\ociram_addr[3]~3_combout ),
	.ociram_addr_4(\ociram_addr[4]~4_combout ),
	.ociram_addr_5(\ociram_addr[5]~5_combout ),
	.ociram_addr_6(\ociram_addr[6]~6_combout ),
	.ociram_addr_7(\ociram_addr[7]~7_combout ),
	.ociram_byteenable_0(\ociram_byteenable[0]~0_combout ),
	.ociram_wr_data_1(\ociram_wr_data[1]~1_combout ),
	.ociram_wr_data_2(\ociram_wr_data[2]~2_combout ),
	.ociram_wr_data_22(\ociram_wr_data[22]~3_combout ),
	.ociram_byteenable_2(\ociram_byteenable[2]~1_combout ),
	.ociram_wr_data_23(\ociram_wr_data[23]~4_combout ),
	.ociram_wr_data_24(\ociram_wr_data[24]~5_combout ),
	.ociram_byteenable_3(\ociram_byteenable[3]~2_combout ),
	.ociram_wr_data_25(\ociram_wr_data[25]~6_combout ),
	.ociram_wr_data_26(\ociram_wr_data[26]~7_combout ),
	.ociram_wr_data_4(\ociram_wr_data[4]~8_combout ),
	.ociram_wr_data_3(\ociram_wr_data[3]~9_combout ),
	.ociram_wr_data_5(\ociram_wr_data[5]~10_combout ),
	.ociram_wr_data_14(\ociram_wr_data[14]~11_combout ),
	.ociram_byteenable_1(\ociram_byteenable[1]~3_combout ),
	.ociram_wr_data_15(\ociram_wr_data[15]~12_combout ),
	.ociram_wr_data_11(\ociram_wr_data[11]~13_combout ),
	.ociram_wr_data_13(\ociram_wr_data[13]~14_combout ),
	.ociram_wr_data_16(\ociram_wr_data[16]~15_combout ),
	.ociram_wr_data_12(\ociram_wr_data[12]~16_combout ),
	.ociram_wr_data_10(\ociram_wr_data[10]~17_combout ),
	.ociram_wr_data_9(\ociram_wr_data[9]~18_combout ),
	.ociram_wr_data_8(\ociram_wr_data[8]~19_combout ),
	.ociram_wr_data_7(\ociram_wr_data[7]~20_combout ),
	.ociram_wr_data_6(\ociram_wr_data[6]~21_combout ),
	.ociram_wr_data_21(\ociram_wr_data[21]~22_combout ),
	.ociram_wr_data_20(\ociram_wr_data[20]~23_combout ),
	.ociram_wr_data_19(\ociram_wr_data[19]~24_combout ),
	.ociram_wr_data_18(\ociram_wr_data[18]~25_combout ),
	.ociram_wr_data_17(\ociram_wr_data[17]~26_combout ),
	.ociram_wr_data_27(\ociram_wr_data[27]~27_combout ),
	.ociram_wr_data_28(\ociram_wr_data[28]~28_combout ),
	.ociram_wr_data_29(\ociram_wr_data[29]~29_combout ),
	.ociram_wr_data_30(\ociram_wr_data[30]~30_combout ),
	.ociram_wr_data_31(\ociram_wr_data[31]~31_combout ),
	.clk_clk(clk_clk));

cyclone10lp_lcell_comb \ociram_wr_en~0 (
	.dataa(write),
	.datab(debugaccess),
	.datac(address_8),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_en~0_combout ),
	.cout());
defparam \ociram_wr_en~0 .lut_mask = 16'hEFFF;
defparam \ociram_wr_en~0 .sum_lutc_input = "datac";

dffeas jtag_ram_wr(
	.clk(clk_clk),
	.d(\jtag_ram_wr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_wr~q ),
	.prn(vcc));
defparam jtag_ram_wr.is_wysiwyg = "true";
defparam jtag_ram_wr.power_up = "low";

cyclone10lp_lcell_comb \ociram_wr_en~1 (
	.dataa(\ociram_wr_en~0_combout ),
	.datab(\jtag_ram_access~q ),
	.datac(\jtag_ram_wr~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ociram_wr_en~1_combout ),
	.cout());
defparam \ociram_wr_en~1 .lut_mask = 16'hFEFE;
defparam \ociram_wr_en~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb ociram_reset_req(
	.dataa(r_early_rst),
	.datab(gnd),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_reset_req~combout ),
	.cout());
defparam ociram_reset_req.lut_mask = 16'hFF55;
defparam ociram_reset_req.sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[0]~0 (
	.dataa(MonDReg_0),
	.datab(writedata_0),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[0]~0_combout ),
	.cout());
defparam \ociram_wr_data[0]~0 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_addr[0]~0 (
	.dataa(\MonAReg[2]~q ),
	.datab(address_0),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[0]~0_combout ),
	.cout());
defparam \ociram_addr[0]~0 .lut_mask = 16'hAACC;
defparam \ociram_addr[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_addr[1]~1 (
	.dataa(\MonAReg[3]~q ),
	.datab(address_1),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[1]~1_combout ),
	.cout());
defparam \ociram_addr[1]~1 .lut_mask = 16'hAACC;
defparam \ociram_addr[1]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_addr[2]~2 (
	.dataa(\MonAReg[4]~q ),
	.datab(address_2),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[2]~2_combout ),
	.cout());
defparam \ociram_addr[2]~2 .lut_mask = 16'hAACC;
defparam \ociram_addr[2]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_addr[3]~3 (
	.dataa(\MonAReg[5]~q ),
	.datab(address_3),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[3]~3_combout ),
	.cout());
defparam \ociram_addr[3]~3 .lut_mask = 16'hAACC;
defparam \ociram_addr[3]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_addr[4]~4 (
	.dataa(\MonAReg[6]~q ),
	.datab(address_4),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[4]~4_combout ),
	.cout());
defparam \ociram_addr[4]~4 .lut_mask = 16'hAACC;
defparam \ociram_addr[4]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_addr[5]~5 (
	.dataa(\MonAReg[7]~q ),
	.datab(address_5),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[5]~5_combout ),
	.cout());
defparam \ociram_addr[5]~5 .lut_mask = 16'hAACC;
defparam \ociram_addr[5]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_addr[6]~6 (
	.dataa(\MonAReg[8]~q ),
	.datab(address_6),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[6]~6_combout ),
	.cout());
defparam \ociram_addr[6]~6 .lut_mask = 16'hAACC;
defparam \ociram_addr[6]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_addr[7]~7 (
	.dataa(\MonAReg[9]~q ),
	.datab(address_7),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[7]~7_combout ),
	.cout());
defparam \ociram_addr[7]~7 .lut_mask = 16'hAACC;
defparam \ociram_addr[7]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_byteenable[0]~0 (
	.dataa(\jtag_ram_access~q ),
	.datab(byteenable_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ociram_byteenable[0]~0_combout ),
	.cout());
defparam \ociram_byteenable[0]~0 .lut_mask = 16'hEEEE;
defparam \ociram_byteenable[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[1]~1 (
	.dataa(MonDReg_1),
	.datab(writedata_1),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[1]~1_combout ),
	.cout());
defparam \ociram_wr_data[1]~1 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[1]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \jtag_ram_wr~0 (
	.dataa(take_action_ocimem_a),
	.datab(\jtag_ram_wr~q ),
	.datac(jdo_35),
	.datad(\MonARegAddrInc[8]~16_combout ),
	.cin(gnd),
	.combout(\jtag_ram_wr~0_combout ),
	.cout());
defparam \jtag_ram_wr~0 .lut_mask = 16'hACFF;
defparam \jtag_ram_wr~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[2]~2 (
	.dataa(MonDReg_2),
	.datab(writedata_2),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[2]~2_combout ),
	.cout());
defparam \ociram_wr_data[2]~2 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[2]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[22]~3 (
	.dataa(MonDReg_22),
	.datab(writedata_22),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[22]~3_combout ),
	.cout());
defparam \ociram_wr_data[22]~3 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[22]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_byteenable[2]~1 (
	.dataa(\jtag_ram_access~q ),
	.datab(byteenable_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ociram_byteenable[2]~1_combout ),
	.cout());
defparam \ociram_byteenable[2]~1 .lut_mask = 16'hEEEE;
defparam \ociram_byteenable[2]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[23]~4 (
	.dataa(MonDReg_23),
	.datab(writedata_23),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[23]~4_combout ),
	.cout());
defparam \ociram_wr_data[23]~4 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[23]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[24]~5 (
	.dataa(MonDReg_24),
	.datab(writedata_24),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[24]~5_combout ),
	.cout());
defparam \ociram_wr_data[24]~5 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[24]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_byteenable[3]~2 (
	.dataa(\jtag_ram_access~q ),
	.datab(byteenable_3),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ociram_byteenable[3]~2_combout ),
	.cout());
defparam \ociram_byteenable[3]~2 .lut_mask = 16'hEEEE;
defparam \ociram_byteenable[3]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[25]~6 (
	.dataa(MonDReg_25),
	.datab(writedata_25),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[25]~6_combout ),
	.cout());
defparam \ociram_wr_data[25]~6 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[25]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[26]~7 (
	.dataa(MonDReg_26),
	.datab(writedata_26),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[26]~7_combout ),
	.cout());
defparam \ociram_wr_data[26]~7 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[26]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[4]~8 (
	.dataa(MonDReg_4),
	.datab(writedata_4),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[4]~8_combout ),
	.cout());
defparam \ociram_wr_data[4]~8 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[4]~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[3]~9 (
	.dataa(MonDReg_3),
	.datab(writedata_3),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[3]~9_combout ),
	.cout());
defparam \ociram_wr_data[3]~9 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[3]~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[5]~10 (
	.dataa(MonDReg_5),
	.datab(writedata_5),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[5]~10_combout ),
	.cout());
defparam \ociram_wr_data[5]~10 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[5]~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[14]~11 (
	.dataa(MonDReg_14),
	.datab(writedata_14),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[14]~11_combout ),
	.cout());
defparam \ociram_wr_data[14]~11 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[14]~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_byteenable[1]~3 (
	.dataa(\jtag_ram_access~q ),
	.datab(byteenable_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ociram_byteenable[1]~3_combout ),
	.cout());
defparam \ociram_byteenable[1]~3 .lut_mask = 16'hEEEE;
defparam \ociram_byteenable[1]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[15]~12 (
	.dataa(MonDReg_15),
	.datab(writedata_15),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[15]~12_combout ),
	.cout());
defparam \ociram_wr_data[15]~12 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[15]~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[11]~13 (
	.dataa(MonDReg_11),
	.datab(writedata_11),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[11]~13_combout ),
	.cout());
defparam \ociram_wr_data[11]~13 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[11]~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[13]~14 (
	.dataa(MonDReg_13),
	.datab(writedata_13),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[13]~14_combout ),
	.cout());
defparam \ociram_wr_data[13]~14 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[13]~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[16]~15 (
	.dataa(MonDReg_16),
	.datab(writedata_16),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[16]~15_combout ),
	.cout());
defparam \ociram_wr_data[16]~15 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[16]~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[12]~16 (
	.dataa(MonDReg_12),
	.datab(writedata_12),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[12]~16_combout ),
	.cout());
defparam \ociram_wr_data[12]~16 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[12]~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[10]~17 (
	.dataa(MonDReg_10),
	.datab(writedata_10),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[10]~17_combout ),
	.cout());
defparam \ociram_wr_data[10]~17 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[10]~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[9]~18 (
	.dataa(MonDReg_9),
	.datab(writedata_9),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[9]~18_combout ),
	.cout());
defparam \ociram_wr_data[9]~18 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[9]~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[8]~19 (
	.dataa(MonDReg_8),
	.datab(writedata_8),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[8]~19_combout ),
	.cout());
defparam \ociram_wr_data[8]~19 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[8]~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[7]~20 (
	.dataa(MonDReg_7),
	.datab(writedata_7),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[7]~20_combout ),
	.cout());
defparam \ociram_wr_data[7]~20 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[7]~20 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[6]~21 (
	.dataa(MonDReg_6),
	.datab(writedata_6),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[6]~21_combout ),
	.cout());
defparam \ociram_wr_data[6]~21 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[6]~21 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[21]~22 (
	.dataa(MonDReg_21),
	.datab(writedata_21),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[21]~22_combout ),
	.cout());
defparam \ociram_wr_data[21]~22 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[21]~22 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[20]~23 (
	.dataa(MonDReg_20),
	.datab(writedata_20),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[20]~23_combout ),
	.cout());
defparam \ociram_wr_data[20]~23 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[20]~23 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[19]~24 (
	.dataa(MonDReg_19),
	.datab(writedata_19),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[19]~24_combout ),
	.cout());
defparam \ociram_wr_data[19]~24 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[19]~24 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[18]~25 (
	.dataa(MonDReg_18),
	.datab(writedata_18),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[18]~25_combout ),
	.cout());
defparam \ociram_wr_data[18]~25 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[18]~25 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[17]~26 (
	.dataa(MonDReg_17),
	.datab(writedata_17),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[17]~26_combout ),
	.cout());
defparam \ociram_wr_data[17]~26 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[17]~26 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[27]~27 (
	.dataa(MonDReg_27),
	.datab(writedata_27),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[27]~27_combout ),
	.cout());
defparam \ociram_wr_data[27]~27 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[27]~27 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[28]~28 (
	.dataa(MonDReg_28),
	.datab(writedata_28),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[28]~28_combout ),
	.cout());
defparam \ociram_wr_data[28]~28 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[28]~28 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[29]~29 (
	.dataa(MonDReg_29),
	.datab(writedata_29),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[29]~29_combout ),
	.cout());
defparam \ociram_wr_data[29]~29 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[29]~29 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[30]~30 (
	.dataa(MonDReg_30),
	.datab(writedata_30),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[30]~30_combout ),
	.cout());
defparam \ociram_wr_data[30]~30 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[30]~30 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ociram_wr_data[31]~31 (
	.dataa(MonDReg_31),
	.datab(writedata_31),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[31]~31_combout ),
	.cout());
defparam \ociram_wr_data[31]~31 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[31]~31 .sum_lutc_input = "datac";

dffeas \MonDReg[0] (
	.clk(clk_clk),
	.d(\MonDReg[0]~0_combout ),
	.asdata(jdo_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~8_combout ),
	.q(MonDReg_0),
	.prn(vcc));
defparam \MonDReg[0] .is_wysiwyg = "true";
defparam \MonDReg[0] .power_up = "low";

dffeas \MonDReg[4] (
	.clk(clk_clk),
	.d(\MonDReg[4]~1_combout ),
	.asdata(jdo_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~8_combout ),
	.q(MonDReg_4),
	.prn(vcc));
defparam \MonDReg[4] .is_wysiwyg = "true";
defparam \MonDReg[4] .power_up = "low";

dffeas \MonDReg[29] (
	.clk(clk_clk),
	.d(\MonDReg[29]~7_combout ),
	.asdata(jdo_32),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~8_combout ),
	.q(MonDReg_29),
	.prn(vcc));
defparam \MonDReg[29] .is_wysiwyg = "true";
defparam \MonDReg[29] .power_up = "low";

dffeas \MonDReg[5] (
	.clk(clk_clk),
	.d(\MonDReg[5]~2_combout ),
	.asdata(jdo_8),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~8_combout ),
	.q(MonDReg_5),
	.prn(vcc));
defparam \MonDReg[5] .is_wysiwyg = "true";
defparam \MonDReg[5] .power_up = "low";

dffeas \MonDReg[15] (
	.clk(clk_clk),
	.d(\MonDReg[15]~3_combout ),
	.asdata(jdo_18),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[15]~26_combout ),
	.q(MonDReg_15),
	.prn(vcc));
defparam \MonDReg[15] .is_wysiwyg = "true";
defparam \MonDReg[15] .power_up = "low";

dffeas \MonDReg[12] (
	.clk(clk_clk),
	.d(\MonDReg[12]~4_combout ),
	.asdata(jdo_15),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~8_combout ),
	.q(MonDReg_12),
	.prn(vcc));
defparam \MonDReg[12] .is_wysiwyg = "true";
defparam \MonDReg[12] .power_up = "low";

dffeas \MonDReg[8] (
	.clk(clk_clk),
	.d(\MonDReg[8]~6_combout ),
	.asdata(jdo_11),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[15]~26_combout ),
	.q(MonDReg_8),
	.prn(vcc));
defparam \MonDReg[8] .is_wysiwyg = "true";
defparam \MonDReg[8] .power_up = "low";

dffeas \MonDReg[18] (
	.clk(clk_clk),
	.d(\MonDReg[18]~5_combout ),
	.asdata(jdo_21),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~8_combout ),
	.q(MonDReg_18),
	.prn(vcc));
defparam \MonDReg[18] .is_wysiwyg = "true";
defparam \MonDReg[18] .power_up = "low";

dffeas waitrequest(
	.clk(clk_clk),
	.d(\waitrequest~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(waitrequest1),
	.prn(vcc));
defparam waitrequest.is_wysiwyg = "true";
defparam waitrequest.power_up = "low";

dffeas \MonDReg[1] (
	.clk(clk_clk),
	.d(\MonDReg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~8_combout ),
	.q(MonDReg_1),
	.prn(vcc));
defparam \MonDReg[1] .is_wysiwyg = "true";
defparam \MonDReg[1] .power_up = "low";

dffeas \MonDReg[2] (
	.clk(clk_clk),
	.d(\MonDReg~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~8_combout ),
	.q(MonDReg_2),
	.prn(vcc));
defparam \MonDReg[2] .is_wysiwyg = "true";
defparam \MonDReg[2] .power_up = "low";

dffeas \MonDReg[3] (
	.clk(clk_clk),
	.d(\MonDReg~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~8_combout ),
	.q(MonDReg_3),
	.prn(vcc));
defparam \MonDReg[3] .is_wysiwyg = "true";
defparam \MonDReg[3] .power_up = "low";

dffeas \MonDReg[16] (
	.clk(clk_clk),
	.d(\MonDReg~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~8_combout ),
	.q(MonDReg_16),
	.prn(vcc));
defparam \MonDReg[16] .is_wysiwyg = "true";
defparam \MonDReg[16] .power_up = "low";

dffeas \MonDReg[25] (
	.clk(clk_clk),
	.d(\MonDReg~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~8_combout ),
	.q(MonDReg_25),
	.prn(vcc));
defparam \MonDReg[25] .is_wysiwyg = "true";
defparam \MonDReg[25] .power_up = "low";

dffeas \MonDReg[27] (
	.clk(clk_clk),
	.d(\MonDReg~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~8_combout ),
	.q(MonDReg_27),
	.prn(vcc));
defparam \MonDReg[27] .is_wysiwyg = "true";
defparam \MonDReg[27] .power_up = "low";

dffeas \MonDReg[26] (
	.clk(clk_clk),
	.d(\MonDReg~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~8_combout ),
	.q(MonDReg_26),
	.prn(vcc));
defparam \MonDReg[26] .is_wysiwyg = "true";
defparam \MonDReg[26] .power_up = "low";

dffeas \MonDReg[24] (
	.clk(clk_clk),
	.d(\MonDReg~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~8_combout ),
	.q(MonDReg_24),
	.prn(vcc));
defparam \MonDReg[24] .is_wysiwyg = "true";
defparam \MonDReg[24] .power_up = "low";

dffeas \MonDReg[20] (
	.clk(clk_clk),
	.d(\MonDReg~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~8_combout ),
	.q(MonDReg_20),
	.prn(vcc));
defparam \MonDReg[20] .is_wysiwyg = "true";
defparam \MonDReg[20] .power_up = "low";

dffeas \MonDReg[19] (
	.clk(clk_clk),
	.d(\MonDReg~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~8_combout ),
	.q(MonDReg_19),
	.prn(vcc));
defparam \MonDReg[19] .is_wysiwyg = "true";
defparam \MonDReg[19] .power_up = "low";

dffeas \MonDReg[22] (
	.clk(clk_clk),
	.d(\MonDReg~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~8_combout ),
	.q(MonDReg_22),
	.prn(vcc));
defparam \MonDReg[22] .is_wysiwyg = "true";
defparam \MonDReg[22] .power_up = "low";

dffeas \MonDReg[23] (
	.clk(clk_clk),
	.d(\MonDReg~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~8_combout ),
	.q(MonDReg_23),
	.prn(vcc));
defparam \MonDReg[23] .is_wysiwyg = "true";
defparam \MonDReg[23] .power_up = "low";

dffeas \MonDReg[17] (
	.clk(clk_clk),
	.d(\MonDReg~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~8_combout ),
	.q(MonDReg_17),
	.prn(vcc));
defparam \MonDReg[17] .is_wysiwyg = "true";
defparam \MonDReg[17] .power_up = "low";

dffeas \MonDReg[31] (
	.clk(clk_clk),
	.d(\MonDReg~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~8_combout ),
	.q(MonDReg_31),
	.prn(vcc));
defparam \MonDReg[31] .is_wysiwyg = "true";
defparam \MonDReg[31] .power_up = "low";

dffeas \MonDReg[30] (
	.clk(clk_clk),
	.d(\MonDReg~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~8_combout ),
	.q(MonDReg_30),
	.prn(vcc));
defparam \MonDReg[30] .is_wysiwyg = "true";
defparam \MonDReg[30] .power_up = "low";

dffeas \MonDReg[28] (
	.clk(clk_clk),
	.d(\MonDReg~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~8_combout ),
	.q(MonDReg_28),
	.prn(vcc));
defparam \MonDReg[28] .is_wysiwyg = "true";
defparam \MonDReg[28] .power_up = "low";

dffeas \MonDReg[14] (
	.clk(clk_clk),
	.d(\MonDReg~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~8_combout ),
	.q(MonDReg_14),
	.prn(vcc));
defparam \MonDReg[14] .is_wysiwyg = "true";
defparam \MonDReg[14] .power_up = "low";

dffeas \MonDReg[11] (
	.clk(clk_clk),
	.d(\MonDReg~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~8_combout ),
	.q(MonDReg_11),
	.prn(vcc));
defparam \MonDReg[11] .is_wysiwyg = "true";
defparam \MonDReg[11] .power_up = "low";

dffeas \MonDReg[13] (
	.clk(clk_clk),
	.d(\MonDReg~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~8_combout ),
	.q(MonDReg_13),
	.prn(vcc));
defparam \MonDReg[13] .is_wysiwyg = "true";
defparam \MonDReg[13] .power_up = "low";

dffeas \MonDReg[10] (
	.clk(clk_clk),
	.d(\MonDReg~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~8_combout ),
	.q(MonDReg_10),
	.prn(vcc));
defparam \MonDReg[10] .is_wysiwyg = "true";
defparam \MonDReg[10] .power_up = "low";

dffeas \MonDReg[9] (
	.clk(clk_clk),
	.d(\MonDReg~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~8_combout ),
	.q(MonDReg_9),
	.prn(vcc));
defparam \MonDReg[9] .is_wysiwyg = "true";
defparam \MonDReg[9] .power_up = "low";

dffeas \MonDReg[7] (
	.clk(clk_clk),
	.d(\MonDReg~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~8_combout ),
	.q(MonDReg_7),
	.prn(vcc));
defparam \MonDReg[7] .is_wysiwyg = "true";
defparam \MonDReg[7] .power_up = "low";

dffeas \MonDReg[6] (
	.clk(clk_clk),
	.d(\MonDReg~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~8_combout ),
	.q(MonDReg_6),
	.prn(vcc));
defparam \MonDReg[6] .is_wysiwyg = "true";
defparam \MonDReg[6] .power_up = "low";

dffeas \MonDReg[21] (
	.clk(clk_clk),
	.d(\MonDReg~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~8_combout ),
	.q(MonDReg_21),
	.prn(vcc));
defparam \MonDReg[21] .is_wysiwyg = "true";
defparam \MonDReg[21] .power_up = "low";

cyclone10lp_lcell_comb \MonARegAddrInc[0]~0 (
	.dataa(\MonAReg[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\MonARegAddrInc[0]~0_combout ),
	.cout(\MonARegAddrInc[0]~1 ));
defparam \MonARegAddrInc[0]~0 .lut_mask = 16'h55AA;
defparam \MonARegAddrInc[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonAReg~0 (
	.dataa(jdo_26),
	.datab(\MonARegAddrInc[0]~0_combout ),
	.datac(take_action_ocimem_a1),
	.datad(jdo_34),
	.cin(gnd),
	.combout(\MonAReg~0_combout ),
	.cout());
defparam \MonAReg~0 .lut_mask = 16'hEFFE;
defparam \MonAReg~0 .sum_lutc_input = "datac";

dffeas \MonAReg[2] (
	.clk(clk_clk),
	.d(\MonAReg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[2]~q ),
	.prn(vcc));
defparam \MonAReg[2] .is_wysiwyg = "true";
defparam \MonAReg[2] .power_up = "low";

cyclone10lp_lcell_comb \MonARegAddrInc[1]~2 (
	.dataa(\MonAReg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[0]~1 ),
	.combout(\MonARegAddrInc[1]~2_combout ),
	.cout(\MonARegAddrInc[1]~3 ));
defparam \MonARegAddrInc[1]~2 .lut_mask = 16'h5A5F;
defparam \MonARegAddrInc[1]~2 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \MonAReg~2 (
	.dataa(jdo_27),
	.datab(\MonARegAddrInc[1]~2_combout ),
	.datac(take_action_ocimem_a1),
	.datad(jdo_34),
	.cin(gnd),
	.combout(\MonAReg~2_combout ),
	.cout());
defparam \MonAReg~2 .lut_mask = 16'hEFFE;
defparam \MonAReg~2 .sum_lutc_input = "datac";

dffeas \MonAReg[3] (
	.clk(clk_clk),
	.d(\MonAReg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[3]~q ),
	.prn(vcc));
defparam \MonAReg[3] .is_wysiwyg = "true";
defparam \MonAReg[3] .power_up = "low";

cyclone10lp_lcell_comb \MonARegAddrInc[2]~4 (
	.dataa(\MonAReg[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[1]~3 ),
	.combout(\MonARegAddrInc[2]~4_combout ),
	.cout(\MonARegAddrInc[2]~5 ));
defparam \MonARegAddrInc[2]~4 .lut_mask = 16'h5AAF;
defparam \MonARegAddrInc[2]~4 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \MonAReg~1 (
	.dataa(jdo_28),
	.datab(\MonARegAddrInc[2]~4_combout ),
	.datac(take_action_ocimem_a1),
	.datad(jdo_34),
	.cin(gnd),
	.combout(\MonAReg~1_combout ),
	.cout());
defparam \MonAReg~1 .lut_mask = 16'hEFFE;
defparam \MonAReg~1 .sum_lutc_input = "datac";

dffeas \MonAReg[4] (
	.clk(clk_clk),
	.d(\MonAReg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[4]~q ),
	.prn(vcc));
defparam \MonAReg[4] .is_wysiwyg = "true";
defparam \MonAReg[4] .power_up = "low";

cyclone10lp_lcell_comb \Equal0~0 (
	.dataa(\MonAReg[2]~q ),
	.datab(gnd),
	.datac(\MonAReg[4]~q ),
	.datad(\MonAReg[3]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hAFFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \jtag_ram_access~0 (
	.dataa(jdo_17),
	.datab(\MonARegAddrInc[8]~16_combout ),
	.datac(take_action_ocimem_a1),
	.datad(jdo_34),
	.cin(gnd),
	.combout(\jtag_ram_access~0_combout ),
	.cout());
defparam \jtag_ram_access~0 .lut_mask = 16'hEFFE;
defparam \jtag_ram_access~0 .sum_lutc_input = "datac";

dffeas \MonAReg[10] (
	.clk(clk_clk),
	.d(\jtag_ram_access~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[10]~q ),
	.prn(vcc));
defparam \MonAReg[10] .is_wysiwyg = "true";
defparam \MonAReg[10] .power_up = "low";

cyclone10lp_lcell_comb \MonARegAddrInc[3]~6 (
	.dataa(\MonAReg[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[2]~5 ),
	.combout(\MonARegAddrInc[3]~6_combout ),
	.cout(\MonARegAddrInc[3]~7 ));
defparam \MonARegAddrInc[3]~6 .lut_mask = 16'h5A5F;
defparam \MonARegAddrInc[3]~6 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \MonAReg~7 (
	.dataa(jdo_29),
	.datab(\MonARegAddrInc[3]~6_combout ),
	.datac(take_action_ocimem_a1),
	.datad(jdo_34),
	.cin(gnd),
	.combout(\MonAReg~7_combout ),
	.cout());
defparam \MonAReg~7 .lut_mask = 16'hEFFE;
defparam \MonAReg~7 .sum_lutc_input = "datac";

dffeas \MonAReg[5] (
	.clk(clk_clk),
	.d(\MonAReg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[5]~q ),
	.prn(vcc));
defparam \MonAReg[5] .is_wysiwyg = "true";
defparam \MonAReg[5] .power_up = "low";

cyclone10lp_lcell_comb \MonARegAddrInc[4]~8 (
	.dataa(\MonAReg[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[3]~7 ),
	.combout(\MonARegAddrInc[4]~8_combout ),
	.cout(\MonARegAddrInc[4]~9 ));
defparam \MonARegAddrInc[4]~8 .lut_mask = 16'h5AAF;
defparam \MonARegAddrInc[4]~8 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \MonAReg~6 (
	.dataa(jdo_30),
	.datab(\MonARegAddrInc[4]~8_combout ),
	.datac(take_action_ocimem_a1),
	.datad(jdo_34),
	.cin(gnd),
	.combout(\MonAReg~6_combout ),
	.cout());
defparam \MonAReg~6 .lut_mask = 16'hEFFE;
defparam \MonAReg~6 .sum_lutc_input = "datac";

dffeas \MonAReg[6] (
	.clk(clk_clk),
	.d(\MonAReg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[6]~q ),
	.prn(vcc));
defparam \MonAReg[6] .is_wysiwyg = "true";
defparam \MonAReg[6] .power_up = "low";

cyclone10lp_lcell_comb \MonARegAddrInc[5]~10 (
	.dataa(\MonAReg[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[4]~9 ),
	.combout(\MonARegAddrInc[5]~10_combout ),
	.cout(\MonARegAddrInc[5]~11 ));
defparam \MonARegAddrInc[5]~10 .lut_mask = 16'h5A5F;
defparam \MonARegAddrInc[5]~10 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \MonAReg~5 (
	.dataa(jdo_31),
	.datab(\MonARegAddrInc[5]~10_combout ),
	.datac(take_action_ocimem_a1),
	.datad(jdo_34),
	.cin(gnd),
	.combout(\MonAReg~5_combout ),
	.cout());
defparam \MonAReg~5 .lut_mask = 16'hEFFE;
defparam \MonAReg~5 .sum_lutc_input = "datac";

dffeas \MonAReg[7] (
	.clk(clk_clk),
	.d(\MonAReg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[7]~q ),
	.prn(vcc));
defparam \MonAReg[7] .is_wysiwyg = "true";
defparam \MonAReg[7] .power_up = "low";

cyclone10lp_lcell_comb \MonARegAddrInc[6]~12 (
	.dataa(\MonAReg[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[5]~11 ),
	.combout(\MonARegAddrInc[6]~12_combout ),
	.cout(\MonARegAddrInc[6]~13 ));
defparam \MonARegAddrInc[6]~12 .lut_mask = 16'h5AAF;
defparam \MonARegAddrInc[6]~12 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \MonAReg~4 (
	.dataa(jdo_32),
	.datab(\MonARegAddrInc[6]~12_combout ),
	.datac(take_action_ocimem_a1),
	.datad(jdo_34),
	.cin(gnd),
	.combout(\MonAReg~4_combout ),
	.cout());
defparam \MonAReg~4 .lut_mask = 16'hEFFE;
defparam \MonAReg~4 .sum_lutc_input = "datac";

dffeas \MonAReg[8] (
	.clk(clk_clk),
	.d(\MonAReg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[8]~q ),
	.prn(vcc));
defparam \MonAReg[8] .is_wysiwyg = "true";
defparam \MonAReg[8] .power_up = "low";

cyclone10lp_lcell_comb \MonARegAddrInc[7]~14 (
	.dataa(\MonAReg[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[6]~13 ),
	.combout(\MonARegAddrInc[7]~14_combout ),
	.cout(\MonARegAddrInc[7]~15 ));
defparam \MonARegAddrInc[7]~14 .lut_mask = 16'h5A5F;
defparam \MonARegAddrInc[7]~14 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \MonAReg~3 (
	.dataa(jdo_33),
	.datab(\MonARegAddrInc[7]~14_combout ),
	.datac(take_action_ocimem_a1),
	.datad(jdo_34),
	.cin(gnd),
	.combout(\MonAReg~3_combout ),
	.cout());
defparam \MonAReg~3 .lut_mask = 16'hEFFE;
defparam \MonAReg~3 .sum_lutc_input = "datac";

dffeas \MonAReg[9] (
	.clk(clk_clk),
	.d(\MonAReg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[9]~q ),
	.prn(vcc));
defparam \MonAReg[9] .is_wysiwyg = "true";
defparam \MonAReg[9] .power_up = "low";

cyclone10lp_lcell_comb \MonARegAddrInc[8]~16 (
	.dataa(\MonAReg[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\MonARegAddrInc[7]~15 ),
	.combout(\MonARegAddrInc[8]~16_combout ),
	.cout());
defparam \MonARegAddrInc[8]~16 .lut_mask = 16'h5A5A;
defparam \MonARegAddrInc[8]~16 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \jtag_ram_rd~0 (
	.dataa(take_action_ocimem_a1),
	.datab(jdo_34),
	.datac(\MonARegAddrInc[8]~16_combout ),
	.datad(jdo_17),
	.cin(gnd),
	.combout(\jtag_ram_rd~0_combout ),
	.cout());
defparam \jtag_ram_rd~0 .lut_mask = 16'h8BFF;
defparam \jtag_ram_rd~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \jtag_ram_rd~1 (
	.dataa(\jtag_ram_rd~0_combout ),
	.datab(take_action_ocimem_b),
	.datac(\jtag_ram_rd~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\jtag_ram_rd~1_combout ),
	.cout());
defparam \jtag_ram_rd~1 .lut_mask = 16'hFEFE;
defparam \jtag_ram_rd~1 .sum_lutc_input = "datac";

dffeas jtag_ram_rd(
	.clk(clk_clk),
	.d(\jtag_ram_rd~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_rd~q ),
	.prn(vcc));
defparam jtag_ram_rd.is_wysiwyg = "true";
defparam jtag_ram_rd.power_up = "low";

dffeas jtag_ram_rd_d1(
	.clk(clk_clk),
	.d(\jtag_ram_rd~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_rd_d1~q ),
	.prn(vcc));
defparam jtag_ram_rd_d1.is_wysiwyg = "true";
defparam jtag_ram_rd_d1.power_up = "low";

cyclone10lp_lcell_comb \MonDReg[0]~0 (
	.dataa(\Equal0~0_combout ),
	.datab(q_a_0),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[0]~0_combout ),
	.cout());
defparam \MonDReg[0]~0 .lut_mask = 16'hAACC;
defparam \MonDReg[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \jtag_rd~0 (
	.dataa(take_action_ocimem_a),
	.datab(\jtag_rd~q ),
	.datac(gnd),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\jtag_rd~0_combout ),
	.cout());
defparam \jtag_rd~0 .lut_mask = 16'hEEFF;
defparam \jtag_rd~0 .sum_lutc_input = "datac";

dffeas jtag_rd(
	.clk(clk_clk),
	.d(\jtag_rd~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_rd~q ),
	.prn(vcc));
defparam jtag_rd.is_wysiwyg = "true";
defparam jtag_rd.power_up = "low";

dffeas jtag_rd_d1(
	.clk(clk_clk),
	.d(\jtag_rd~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_rd_d1~q ),
	.prn(vcc));
defparam jtag_rd_d1.is_wysiwyg = "true";
defparam jtag_rd_d1.power_up = "low";

cyclone10lp_lcell_comb \MonDReg[0]~8 (
	.dataa(gnd),
	.datab(take_action_ocimem_a),
	.datac(\jtag_rd_d1~q ),
	.datad(jdo_35),
	.cin(gnd),
	.combout(\MonDReg[0]~8_combout ),
	.cout());
defparam \MonDReg[0]~8 .lut_mask = 16'hF3C0;
defparam \MonDReg[0]~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg[4]~1 (
	.dataa(\Equal0~0_combout ),
	.datab(q_a_4),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[4]~1_combout ),
	.cout());
defparam \MonDReg[4]~1 .lut_mask = 16'hAACC;
defparam \MonDReg[4]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal0~1 (
	.dataa(\MonAReg[4]~q ),
	.datab(gnd),
	.datac(\MonAReg[2]~q ),
	.datad(\MonAReg[3]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'hAFFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg[29]~7 (
	.dataa(\Equal0~1_combout ),
	.datab(q_a_29),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[29]~7_combout ),
	.cout());
defparam \MonDReg[29]~7 .lut_mask = 16'hAACC;
defparam \MonDReg[29]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal0~2 (
	.dataa(gnd),
	.datab(\MonAReg[2]~q ),
	.datac(\MonAReg[4]~q ),
	.datad(\MonAReg[3]~q ),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
defparam \Equal0~2 .lut_mask = 16'h3FFF;
defparam \Equal0~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg[5]~2 (
	.dataa(\Equal0~2_combout ),
	.datab(q_a_5),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[5]~2_combout ),
	.cout());
defparam \MonDReg[5]~2 .lut_mask = 16'hAACC;
defparam \MonDReg[5]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \cfgrom_readdata[15]~0 (
	.dataa(\MonAReg[3]~q ),
	.datab(gnd),
	.datac(\MonAReg[2]~q ),
	.datad(\MonAReg[4]~q ),
	.cin(gnd),
	.combout(\cfgrom_readdata[15]~0_combout ),
	.cout());
defparam \cfgrom_readdata[15]~0 .lut_mask = 16'hAFFA;
defparam \cfgrom_readdata[15]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg[15]~3 (
	.dataa(\cfgrom_readdata[15]~0_combout ),
	.datab(q_a_15),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[15]~3_combout ),
	.cout());
defparam \MonDReg[15]~3 .lut_mask = 16'hCC55;
defparam \MonDReg[15]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg[15]~26 (
	.dataa(take_action_ocimem_b),
	.datab(\jtag_rd_d1~q ),
	.datac(gnd),
	.datad(take_action_ocimem_a),
	.cin(gnd),
	.combout(\MonDReg[15]~26_combout ),
	.cout());
defparam \MonDReg[15]~26 .lut_mask = 16'hEEFF;
defparam \MonDReg[15]~26 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg[12]~4 (
	.dataa(\Equal0~0_combout ),
	.datab(q_a_12),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[12]~4_combout ),
	.cout());
defparam \MonDReg[12]~4 .lut_mask = 16'hAACC;
defparam \MonDReg[12]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \cfgrom_readdata[8]~1 (
	.dataa(\MonAReg[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\MonAReg[4]~q ),
	.cin(gnd),
	.combout(\cfgrom_readdata[8]~1_combout ),
	.cout());
defparam \cfgrom_readdata[8]~1 .lut_mask = 16'hAAFF;
defparam \cfgrom_readdata[8]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg[8]~6 (
	.dataa(\cfgrom_readdata[8]~1_combout ),
	.datab(q_a_8),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[8]~6_combout ),
	.cout());
defparam \MonDReg[8]~6 .lut_mask = 16'hAACC;
defparam \MonDReg[8]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal0~3 (
	.dataa(\MonAReg[3]~q ),
	.datab(gnd),
	.datac(\MonAReg[2]~q ),
	.datad(\MonAReg[4]~q ),
	.cin(gnd),
	.combout(\Equal0~3_combout ),
	.cout());
defparam \Equal0~3 .lut_mask = 16'hAFFF;
defparam \Equal0~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg[18]~5 (
	.dataa(\Equal0~3_combout ),
	.datab(q_a_18),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[18]~5_combout ),
	.cout());
defparam \MonDReg[18]~5 .lut_mask = 16'hAACC;
defparam \MonDReg[18]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \jtag_ram_access~1 (
	.dataa(\jtag_ram_access~0_combout ),
	.datab(\MonARegAddrInc[8]~16_combout ),
	.datac(take_action_ocimem_b),
	.datad(take_action_ocimem_a1),
	.cin(gnd),
	.combout(\jtag_ram_access~1_combout ),
	.cout());
defparam \jtag_ram_access~1 .lut_mask = 16'hF377;
defparam \jtag_ram_access~1 .sum_lutc_input = "datac";

dffeas jtag_ram_access(
	.clk(clk_clk),
	.d(\jtag_ram_access~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_access~q ),
	.prn(vcc));
defparam jtag_ram_access.is_wysiwyg = "true";
defparam jtag_ram_access.power_up = "low";

cyclone10lp_lcell_comb \waitrequest~0 (
	.dataa(write),
	.datab(\jtag_ram_access~q ),
	.datac(address_8),
	.datad(waitrequest1),
	.cin(gnd),
	.combout(\waitrequest~0_combout ),
	.cout());
defparam \waitrequest~0 .lut_mask = 16'hEFFF;
defparam \waitrequest~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \avalon_ociram_readdata_ready~0 (
	.dataa(read),
	.datab(address_8),
	.datac(\jtag_ram_access~q ),
	.datad(write),
	.cin(gnd),
	.combout(\avalon_ociram_readdata_ready~0_combout ),
	.cout());
defparam \avalon_ociram_readdata_ready~0 .lut_mask = 16'hEFFF;
defparam \avalon_ociram_readdata_ready~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \avalon_ociram_readdata_ready~1 (
	.dataa(waitrequest1),
	.datab(\avalon_ociram_readdata_ready~0_combout ),
	.datac(write),
	.datad(\avalon_ociram_readdata_ready~q ),
	.cin(gnd),
	.combout(\avalon_ociram_readdata_ready~1_combout ),
	.cout());
defparam \avalon_ociram_readdata_ready~1 .lut_mask = 16'hFFFE;
defparam \avalon_ociram_readdata_ready~1 .sum_lutc_input = "datac";

dffeas avalon_ociram_readdata_ready(
	.clk(clk_clk),
	.d(\avalon_ociram_readdata_ready~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\avalon_ociram_readdata_ready~q ),
	.prn(vcc));
defparam avalon_ociram_readdata_ready.is_wysiwyg = "true";
defparam avalon_ociram_readdata_ready.power_up = "low";

cyclone10lp_lcell_comb \waitrequest~1 (
	.dataa(\waitrequest~0_combout ),
	.datab(read),
	.datac(\avalon_ociram_readdata_ready~q ),
	.datad(write),
	.cin(gnd),
	.combout(\waitrequest~1_combout ),
	.cout());
defparam \waitrequest~1 .lut_mask = 16'hBFFF;
defparam \waitrequest~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg~9 (
	.dataa(jdo_4),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_1),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~9_combout ),
	.cout());
defparam \MonDReg~9 .lut_mask = 16'hFAFC;
defparam \MonDReg~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg~10 (
	.dataa(jdo_5),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_2),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~10_combout ),
	.cout());
defparam \MonDReg~10 .lut_mask = 16'hFAFC;
defparam \MonDReg~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg~11 (
	.dataa(jdo_6),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_3),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~11_combout ),
	.cout());
defparam \MonDReg~11 .lut_mask = 16'hFAFC;
defparam \MonDReg~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg~12 (
	.dataa(jdo_19),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_16),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~12_combout ),
	.cout());
defparam \MonDReg~12 .lut_mask = 16'hFAFC;
defparam \MonDReg~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg~13 (
	.dataa(jdo_28),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_25),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~13_combout ),
	.cout());
defparam \MonDReg~13 .lut_mask = 16'hFAFC;
defparam \MonDReg~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg~14 (
	.dataa(jdo_30),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_27),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~14_combout ),
	.cout());
defparam \MonDReg~14 .lut_mask = 16'hFAFC;
defparam \MonDReg~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg~15 (
	.dataa(jdo_29),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_26),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~15_combout ),
	.cout());
defparam \MonDReg~15 .lut_mask = 16'hFAFC;
defparam \MonDReg~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg~16 (
	.dataa(jdo_27),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_24),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~16_combout ),
	.cout());
defparam \MonDReg~16 .lut_mask = 16'hFAFC;
defparam \MonDReg~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg~17 (
	.dataa(jdo_23),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_20),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~17_combout ),
	.cout());
defparam \MonDReg~17 .lut_mask = 16'hFAFC;
defparam \MonDReg~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg~18 (
	.dataa(jdo_22),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_19),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~18_combout ),
	.cout());
defparam \MonDReg~18 .lut_mask = 16'hFAFC;
defparam \MonDReg~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg~19 (
	.dataa(jdo_25),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_22),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~19_combout ),
	.cout());
defparam \MonDReg~19 .lut_mask = 16'hFAFC;
defparam \MonDReg~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg~20 (
	.dataa(jdo_26),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_23),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~20_combout ),
	.cout());
defparam \MonDReg~20 .lut_mask = 16'hFAFC;
defparam \MonDReg~20 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg~21 (
	.dataa(jdo_20),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_17),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~21_combout ),
	.cout());
defparam \MonDReg~21 .lut_mask = 16'hFAFC;
defparam \MonDReg~21 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg~22 (
	.dataa(jdo_34),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_31),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~22_combout ),
	.cout());
defparam \MonDReg~22 .lut_mask = 16'hFAFC;
defparam \MonDReg~22 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg~23 (
	.dataa(jdo_33),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_30),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~23_combout ),
	.cout());
defparam \MonDReg~23 .lut_mask = 16'hFAFC;
defparam \MonDReg~23 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg~24 (
	.dataa(jdo_31),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_28),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~24_combout ),
	.cout());
defparam \MonDReg~24 .lut_mask = 16'hFAFC;
defparam \MonDReg~24 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg~25 (
	.dataa(jdo_17),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_14),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~25_combout ),
	.cout());
defparam \MonDReg~25 .lut_mask = 16'hFAFC;
defparam \MonDReg~25 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg~27 (
	.dataa(jdo_14),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_11),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~27_combout ),
	.cout());
defparam \MonDReg~27 .lut_mask = 16'hFAFC;
defparam \MonDReg~27 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg~28 (
	.dataa(jdo_16),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_13),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~28_combout ),
	.cout());
defparam \MonDReg~28 .lut_mask = 16'hFAFC;
defparam \MonDReg~28 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg~29 (
	.dataa(jdo_13),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_10),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~29_combout ),
	.cout());
defparam \MonDReg~29 .lut_mask = 16'hFAFC;
defparam \MonDReg~29 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg~30 (
	.dataa(jdo_12),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_9),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~30_combout ),
	.cout());
defparam \MonDReg~30 .lut_mask = 16'hFAFC;
defparam \MonDReg~30 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg~31 (
	.dataa(jdo_10),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_7),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~31_combout ),
	.cout());
defparam \MonDReg~31 .lut_mask = 16'hFAFC;
defparam \MonDReg~31 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg~32 (
	.dataa(jdo_9),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_6),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~32_combout ),
	.cout());
defparam \MonDReg~32 .lut_mask = 16'hFAFC;
defparam \MonDReg~32 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MonDReg~33 (
	.dataa(jdo_24),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_21),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~33_combout ),
	.cout());
defparam \MonDReg~33 .lut_mask = 16'hFAFC;
defparam \MonDReg~33 .sum_lutc_input = "datac";

endmodule

module processor_processor_nios2_gen2_0_cpu_ociram_sp_ram_module (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_22,
	q_a_23,
	q_a_24,
	q_a_25,
	q_a_26,
	q_a_4,
	q_a_3,
	q_a_5,
	q_a_14,
	q_a_15,
	q_a_11,
	q_a_13,
	q_a_16,
	q_a_12,
	q_a_10,
	q_a_9,
	q_a_8,
	q_a_7,
	q_a_6,
	q_a_21,
	q_a_20,
	q_a_19,
	q_a_18,
	q_a_17,
	q_a_27,
	q_a_28,
	q_a_29,
	q_a_30,
	q_a_31,
	ociram_wr_en,
	ociram_reset_req,
	ociram_wr_data_0,
	ociram_addr_0,
	ociram_addr_1,
	ociram_addr_2,
	ociram_addr_3,
	ociram_addr_4,
	ociram_addr_5,
	ociram_addr_6,
	ociram_addr_7,
	ociram_byteenable_0,
	ociram_wr_data_1,
	ociram_wr_data_2,
	ociram_wr_data_22,
	ociram_byteenable_2,
	ociram_wr_data_23,
	ociram_wr_data_24,
	ociram_byteenable_3,
	ociram_wr_data_25,
	ociram_wr_data_26,
	ociram_wr_data_4,
	ociram_wr_data_3,
	ociram_wr_data_5,
	ociram_wr_data_14,
	ociram_byteenable_1,
	ociram_wr_data_15,
	ociram_wr_data_11,
	ociram_wr_data_13,
	ociram_wr_data_16,
	ociram_wr_data_12,
	ociram_wr_data_10,
	ociram_wr_data_9,
	ociram_wr_data_8,
	ociram_wr_data_7,
	ociram_wr_data_6,
	ociram_wr_data_21,
	ociram_wr_data_20,
	ociram_wr_data_19,
	ociram_wr_data_18,
	ociram_wr_data_17,
	ociram_wr_data_27,
	ociram_wr_data_28,
	ociram_wr_data_29,
	ociram_wr_data_30,
	ociram_wr_data_31,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_22;
output 	q_a_23;
output 	q_a_24;
output 	q_a_25;
output 	q_a_26;
output 	q_a_4;
output 	q_a_3;
output 	q_a_5;
output 	q_a_14;
output 	q_a_15;
output 	q_a_11;
output 	q_a_13;
output 	q_a_16;
output 	q_a_12;
output 	q_a_10;
output 	q_a_9;
output 	q_a_8;
output 	q_a_7;
output 	q_a_6;
output 	q_a_21;
output 	q_a_20;
output 	q_a_19;
output 	q_a_18;
output 	q_a_17;
output 	q_a_27;
output 	q_a_28;
output 	q_a_29;
output 	q_a_30;
output 	q_a_31;
input 	ociram_wr_en;
input 	ociram_reset_req;
input 	ociram_wr_data_0;
input 	ociram_addr_0;
input 	ociram_addr_1;
input 	ociram_addr_2;
input 	ociram_addr_3;
input 	ociram_addr_4;
input 	ociram_addr_5;
input 	ociram_addr_6;
input 	ociram_addr_7;
input 	ociram_byteenable_0;
input 	ociram_wr_data_1;
input 	ociram_wr_data_2;
input 	ociram_wr_data_22;
input 	ociram_byteenable_2;
input 	ociram_wr_data_23;
input 	ociram_wr_data_24;
input 	ociram_byteenable_3;
input 	ociram_wr_data_25;
input 	ociram_wr_data_26;
input 	ociram_wr_data_4;
input 	ociram_wr_data_3;
input 	ociram_wr_data_5;
input 	ociram_wr_data_14;
input 	ociram_byteenable_1;
input 	ociram_wr_data_15;
input 	ociram_wr_data_11;
input 	ociram_wr_data_13;
input 	ociram_wr_data_16;
input 	ociram_wr_data_12;
input 	ociram_wr_data_10;
input 	ociram_wr_data_9;
input 	ociram_wr_data_8;
input 	ociram_wr_data_7;
input 	ociram_wr_data_6;
input 	ociram_wr_data_21;
input 	ociram_wr_data_20;
input 	ociram_wr_data_19;
input 	ociram_wr_data_18;
input 	ociram_wr_data_17;
input 	ociram_wr_data_27;
input 	ociram_wr_data_28;
input 	ociram_wr_data_29;
input 	ociram_wr_data_30;
input 	ociram_wr_data_31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



processor_altsyncram_1 the_altsyncram(
	.q_a({q_a_31,q_a_30,q_a_29,q_a_28,q_a_27,q_a_26,q_a_25,q_a_24,q_a_23,q_a_22,q_a_21,q_a_20,q_a_19,q_a_18,q_a_17,q_a_16,q_a_15,q_a_14,q_a_13,q_a_12,q_a_11,q_a_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.wren_a(ociram_wr_en),
	.clocken0(ociram_reset_req),
	.data_a({ociram_wr_data_31,ociram_wr_data_30,ociram_wr_data_29,ociram_wr_data_28,ociram_wr_data_27,ociram_wr_data_26,ociram_wr_data_25,ociram_wr_data_24,ociram_wr_data_23,ociram_wr_data_22,ociram_wr_data_21,ociram_wr_data_20,ociram_wr_data_19,ociram_wr_data_18,ociram_wr_data_17,
ociram_wr_data_16,ociram_wr_data_15,ociram_wr_data_14,ociram_wr_data_13,ociram_wr_data_12,ociram_wr_data_11,ociram_wr_data_10,ociram_wr_data_9,ociram_wr_data_8,ociram_wr_data_7,ociram_wr_data_6,ociram_wr_data_5,ociram_wr_data_4,ociram_wr_data_3,ociram_wr_data_2,
ociram_wr_data_1,ociram_wr_data_0}),
	.address_a({gnd,gnd,gnd,gnd,gnd,ociram_addr_7,ociram_addr_6,ociram_addr_5,ociram_addr_4,ociram_addr_3,ociram_addr_2,ociram_addr_1,ociram_addr_0}),
	.byteena_a({ociram_byteenable_3,ociram_byteenable_2,ociram_byteenable_1,ociram_byteenable_0}),
	.clock0(clk_clk));

endmodule

module processor_altsyncram_1 (
	q_a,
	wren_a,
	clocken0,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	wren_a;
input 	clocken0;
input 	[31:0] data_a;
input 	[12:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



processor_altsyncram_3c71 auto_generated(
	.q_a({q_a[31],q_a[30],q_a[29],q_a[28],q_a[27],q_a[26],q_a[25],q_a[24],q_a[23],q_a[22],q_a[21],q_a[20],q_a[19],q_a[18],q_a[17],q_a[16],q_a[15],q_a[14],q_a[13],q_a[12],q_a[11],q_a[10],q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.wren_a(wren_a),
	.clocken0(clocken0),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.byteena_a({byteena_a[3],byteena_a[2],byteena_a[1],byteena_a[0]}),
	.clock0(clock0));

endmodule

module processor_altsyncram_3c71 (
	q_a,
	wren_a,
	clocken0,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	wren_a;
input 	clocken0;
input 	[31:0] data_a;
input 	[7:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;
wire [143:0] ram_block1a24_PORTADATAOUT_bus;
wire [143:0] ram_block1a25_PORTADATAOUT_bus;
wire [143:0] ram_block1a26_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;
wire [143:0] ram_block1a27_PORTADATAOUT_bus;
wire [143:0] ram_block1a28_PORTADATAOUT_bus;
wire [143:0] ram_block1a29_PORTADATAOUT_bus;
wire [143:0] ram_block1a30_PORTADATAOUT_bus;
wire [143:0] ram_block1a31_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[22] = ram_block1a22_PORTADATAOUT_bus[0];

assign q_a[23] = ram_block1a23_PORTADATAOUT_bus[0];

assign q_a[24] = ram_block1a24_PORTADATAOUT_bus[0];

assign q_a[25] = ram_block1a25_PORTADATAOUT_bus[0];

assign q_a[26] = ram_block1a26_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[14] = ram_block1a14_PORTADATAOUT_bus[0];

assign q_a[15] = ram_block1a15_PORTADATAOUT_bus[0];

assign q_a[11] = ram_block1a11_PORTADATAOUT_bus[0];

assign q_a[13] = ram_block1a13_PORTADATAOUT_bus[0];

assign q_a[16] = ram_block1a16_PORTADATAOUT_bus[0];

assign q_a[12] = ram_block1a12_PORTADATAOUT_bus[0];

assign q_a[10] = ram_block1a10_PORTADATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[21] = ram_block1a21_PORTADATAOUT_bus[0];

assign q_a[20] = ram_block1a20_PORTADATAOUT_bus[0];

assign q_a[19] = ram_block1a19_PORTADATAOUT_bus[0];

assign q_a[18] = ram_block1a18_PORTADATAOUT_bus[0];

assign q_a[17] = ram_block1a17_PORTADATAOUT_bus[0];

assign q_a[27] = ram_block1a27_PORTADATAOUT_bus[0];

assign q_a[28] = ram_block1a28_PORTADATAOUT_bus[0];

assign q_a[29] = ram_block1a29_PORTADATAOUT_bus[0];

assign q_a[30] = ram_block1a30_PORTADATAOUT_bus[0];

assign q_a[31] = ram_block1a31_PORTADATAOUT_bus[0];

cyclone10lp_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "single_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 8;
defparam ram_block1a0.port_a_byte_enable_mask_width = 1;
defparam ram_block1a0.port_a_byte_size = 1;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 255;
defparam ram_block1a0.port_a_logical_ram_depth = 256;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "single_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 8;
defparam ram_block1a1.port_a_byte_enable_mask_width = 1;
defparam ram_block1a1.port_a_byte_size = 1;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 255;
defparam ram_block1a1.port_a_logical_ram_depth = 256;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "single_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 8;
defparam ram_block1a2.port_a_byte_enable_mask_width = 1;
defparam ram_block1a2.port_a_byte_size = 1;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 255;
defparam ram_block1a2.port_a_logical_ram_depth = 256;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.operation_mode = "single_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 8;
defparam ram_block1a22.port_a_byte_enable_mask_width = 1;
defparam ram_block1a22.port_a_byte_size = 1;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 255;
defparam ram_block1a22.port_a_logical_ram_depth = 256;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.operation_mode = "single_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 8;
defparam ram_block1a23.port_a_byte_enable_mask_width = 1;
defparam ram_block1a23.port_a_byte_size = 1;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 255;
defparam ram_block1a23.port_a_logical_ram_depth = 256;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a24_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.operation_mode = "single_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 8;
defparam ram_block1a24.port_a_byte_enable_mask_width = 1;
defparam ram_block1a24.port_a_byte_size = 1;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 255;
defparam ram_block1a24.port_a_logical_ram_depth = 256;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a25_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.operation_mode = "single_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 8;
defparam ram_block1a25.port_a_byte_enable_mask_width = 1;
defparam ram_block1a25.port_a_byte_size = 1;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 255;
defparam ram_block1a25.port_a_logical_ram_depth = 256;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a26_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.operation_mode = "single_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 8;
defparam ram_block1a26.port_a_byte_enable_mask_width = 1;
defparam ram_block1a26.port_a_byte_size = 1;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 255;
defparam ram_block1a26.port_a_logical_ram_depth = 256;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "single_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 8;
defparam ram_block1a4.port_a_byte_enable_mask_width = 1;
defparam ram_block1a4.port_a_byte_size = 1;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 255;
defparam ram_block1a4.port_a_logical_ram_depth = 256;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "single_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 8;
defparam ram_block1a3.port_a_byte_enable_mask_width = 1;
defparam ram_block1a3.port_a_byte_size = 1;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 255;
defparam ram_block1a3.port_a_logical_ram_depth = 256;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "single_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 8;
defparam ram_block1a5.port_a_byte_enable_mask_width = 1;
defparam ram_block1a5.port_a_byte_size = 1;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 255;
defparam ram_block1a5.port_a_logical_ram_depth = 256;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.operation_mode = "single_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 8;
defparam ram_block1a14.port_a_byte_enable_mask_width = 1;
defparam ram_block1a14.port_a_byte_size = 1;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 255;
defparam ram_block1a14.port_a_logical_ram_depth = 256;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.operation_mode = "single_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 8;
defparam ram_block1a15.port_a_byte_enable_mask_width = 1;
defparam ram_block1a15.port_a_byte_size = 1;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 255;
defparam ram_block1a15.port_a_logical_ram_depth = 256;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.operation_mode = "single_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 8;
defparam ram_block1a11.port_a_byte_enable_mask_width = 1;
defparam ram_block1a11.port_a_byte_size = 1;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 255;
defparam ram_block1a11.port_a_logical_ram_depth = 256;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.operation_mode = "single_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 8;
defparam ram_block1a13.port_a_byte_enable_mask_width = 1;
defparam ram_block1a13.port_a_byte_size = 1;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 255;
defparam ram_block1a13.port_a_logical_ram_depth = 256;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.operation_mode = "single_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 8;
defparam ram_block1a16.port_a_byte_enable_mask_width = 1;
defparam ram_block1a16.port_a_byte_size = 1;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 255;
defparam ram_block1a16.port_a_logical_ram_depth = 256;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.operation_mode = "single_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 8;
defparam ram_block1a12.port_a_byte_enable_mask_width = 1;
defparam ram_block1a12.port_a_byte_size = 1;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 255;
defparam ram_block1a12.port_a_logical_ram_depth = 256;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.operation_mode = "single_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 8;
defparam ram_block1a10.port_a_byte_enable_mask_width = 1;
defparam ram_block1a10.port_a_byte_size = 1;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 255;
defparam ram_block1a10.port_a_logical_ram_depth = 256;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "single_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 8;
defparam ram_block1a9.port_a_byte_enable_mask_width = 1;
defparam ram_block1a9.port_a_byte_size = 1;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 255;
defparam ram_block1a9.port_a_logical_ram_depth = 256;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "single_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 8;
defparam ram_block1a8.port_a_byte_enable_mask_width = 1;
defparam ram_block1a8.port_a_byte_size = 1;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 255;
defparam ram_block1a8.port_a_logical_ram_depth = 256;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "single_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 8;
defparam ram_block1a7.port_a_byte_enable_mask_width = 1;
defparam ram_block1a7.port_a_byte_size = 1;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 255;
defparam ram_block1a7.port_a_logical_ram_depth = 256;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "single_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 8;
defparam ram_block1a6.port_a_byte_enable_mask_width = 1;
defparam ram_block1a6.port_a_byte_size = 1;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 255;
defparam ram_block1a6.port_a_logical_ram_depth = 256;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.operation_mode = "single_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 8;
defparam ram_block1a21.port_a_byte_enable_mask_width = 1;
defparam ram_block1a21.port_a_byte_size = 1;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 255;
defparam ram_block1a21.port_a_logical_ram_depth = 256;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.operation_mode = "single_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 8;
defparam ram_block1a20.port_a_byte_enable_mask_width = 1;
defparam ram_block1a20.port_a_byte_size = 1;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 255;
defparam ram_block1a20.port_a_logical_ram_depth = 256;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.operation_mode = "single_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 8;
defparam ram_block1a19.port_a_byte_enable_mask_width = 1;
defparam ram_block1a19.port_a_byte_size = 1;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 255;
defparam ram_block1a19.port_a_logical_ram_depth = 256;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.operation_mode = "single_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 8;
defparam ram_block1a18.port_a_byte_enable_mask_width = 1;
defparam ram_block1a18.port_a_byte_size = 1;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 255;
defparam ram_block1a18.port_a_logical_ram_depth = 256;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.operation_mode = "single_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 8;
defparam ram_block1a17.port_a_byte_enable_mask_width = 1;
defparam ram_block1a17.port_a_byte_size = 1;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 255;
defparam ram_block1a17.port_a_logical_ram_depth = 256;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a27_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.operation_mode = "single_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 8;
defparam ram_block1a27.port_a_byte_enable_mask_width = 1;
defparam ram_block1a27.port_a_byte_size = 1;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 255;
defparam ram_block1a27.port_a_logical_ram_depth = 256;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a28_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.operation_mode = "single_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 8;
defparam ram_block1a28.port_a_byte_enable_mask_width = 1;
defparam ram_block1a28.port_a_byte_size = 1;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 255;
defparam ram_block1a28.port_a_logical_ram_depth = 256;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a29_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.operation_mode = "single_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 8;
defparam ram_block1a29.port_a_byte_enable_mask_width = 1;
defparam ram_block1a29.port_a_byte_size = 1;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 255;
defparam ram_block1a29.port_a_logical_ram_depth = 256;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a30_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.operation_mode = "single_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 8;
defparam ram_block1a30.port_a_byte_enable_mask_width = 1;
defparam ram_block1a30.port_a_byte_size = 1;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 255;
defparam ram_block1a30.port_a_logical_ram_depth = 256;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a31_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_nios2_oci:the_processor_nios2_gen2_0_cpu_nios2_oci|processor_nios2_gen2_0_cpu_nios2_ocimem:the_processor_nios2_gen2_0_cpu_nios2_ocimem|processor_nios2_gen2_0_cpu_ociram_sp_ram_module:processor_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_3c71:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.operation_mode = "single_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 8;
defparam ram_block1a31.port_a_byte_enable_mask_width = 1;
defparam ram_block1a31.port_a_byte_size = 1;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 255;
defparam ram_block1a31.port_a_logical_ram_depth = 256;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.ram_block_type = "auto";

endmodule

module processor_processor_nios2_gen2_0_cpu_register_bank_a_module (
	q_b_7,
	q_b_6,
	q_b_5,
	q_b_4,
	q_b_3,
	q_b_2,
	q_b_1,
	q_b_0,
	q_b_16,
	q_b_15,
	q_b_14,
	q_b_13,
	q_b_12,
	q_b_11,
	q_b_10,
	q_b_9,
	q_b_8,
	q_b_31,
	q_b_30,
	q_b_29,
	q_b_28,
	q_b_27,
	q_b_26,
	q_b_25,
	q_b_24,
	q_b_23,
	q_b_22,
	q_b_21,
	q_b_20,
	q_b_19,
	q_b_18,
	q_b_17,
	W_rf_wren,
	W_rf_wr_data_0,
	R_dst_regnum_0,
	R_dst_regnum_1,
	R_dst_regnum_2,
	R_dst_regnum_3,
	R_dst_regnum_4,
	W_rf_wr_data_1,
	W_rf_wr_data_2,
	W_rf_wr_data_3,
	W_rf_wr_data_4,
	W_rf_wr_data_5,
	W_rf_wr_data_6,
	W_rf_wr_data_7,
	D_iw_27,
	D_iw_28,
	D_iw_29,
	D_iw_30,
	D_iw_31,
	W_rf_wr_data_16,
	W_rf_wr_data_15,
	W_rf_wr_data_14,
	W_rf_wr_data_13,
	W_rf_wr_data_12,
	W_rf_wr_data_11,
	W_rf_wr_data_10,
	W_rf_wr_data_9,
	W_rf_wr_data_8,
	W_rf_wr_data_31,
	W_rf_wr_data_30,
	W_rf_wr_data_29,
	W_rf_wr_data_28,
	W_rf_wr_data_27,
	W_rf_wr_data_26,
	W_rf_wr_data_25,
	W_rf_wr_data_24,
	W_rf_wr_data_23,
	W_rf_wr_data_22,
	W_rf_wr_data_21,
	W_rf_wr_data_20,
	W_rf_wr_data_19,
	W_rf_wr_data_18,
	W_rf_wr_data_17,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_7;
output 	q_b_6;
output 	q_b_5;
output 	q_b_4;
output 	q_b_3;
output 	q_b_2;
output 	q_b_1;
output 	q_b_0;
output 	q_b_16;
output 	q_b_15;
output 	q_b_14;
output 	q_b_13;
output 	q_b_12;
output 	q_b_11;
output 	q_b_10;
output 	q_b_9;
output 	q_b_8;
output 	q_b_31;
output 	q_b_30;
output 	q_b_29;
output 	q_b_28;
output 	q_b_27;
output 	q_b_26;
output 	q_b_25;
output 	q_b_24;
output 	q_b_23;
output 	q_b_22;
output 	q_b_21;
output 	q_b_20;
output 	q_b_19;
output 	q_b_18;
output 	q_b_17;
input 	W_rf_wren;
input 	W_rf_wr_data_0;
input 	R_dst_regnum_0;
input 	R_dst_regnum_1;
input 	R_dst_regnum_2;
input 	R_dst_regnum_3;
input 	R_dst_regnum_4;
input 	W_rf_wr_data_1;
input 	W_rf_wr_data_2;
input 	W_rf_wr_data_3;
input 	W_rf_wr_data_4;
input 	W_rf_wr_data_5;
input 	W_rf_wr_data_6;
input 	W_rf_wr_data_7;
input 	D_iw_27;
input 	D_iw_28;
input 	D_iw_29;
input 	D_iw_30;
input 	D_iw_31;
input 	W_rf_wr_data_16;
input 	W_rf_wr_data_15;
input 	W_rf_wr_data_14;
input 	W_rf_wr_data_13;
input 	W_rf_wr_data_12;
input 	W_rf_wr_data_11;
input 	W_rf_wr_data_10;
input 	W_rf_wr_data_9;
input 	W_rf_wr_data_8;
input 	W_rf_wr_data_31;
input 	W_rf_wr_data_30;
input 	W_rf_wr_data_29;
input 	W_rf_wr_data_28;
input 	W_rf_wr_data_27;
input 	W_rf_wr_data_26;
input 	W_rf_wr_data_25;
input 	W_rf_wr_data_24;
input 	W_rf_wr_data_23;
input 	W_rf_wr_data_22;
input 	W_rf_wr_data_21;
input 	W_rf_wr_data_20;
input 	W_rf_wr_data_19;
input 	W_rf_wr_data_18;
input 	W_rf_wr_data_17;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



processor_altsyncram_2 the_altsyncram(
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.wren_a(W_rf_wren),
	.data_a({W_rf_wr_data_31,W_rf_wr_data_30,W_rf_wr_data_29,W_rf_wr_data_28,W_rf_wr_data_27,W_rf_wr_data_26,W_rf_wr_data_25,W_rf_wr_data_24,W_rf_wr_data_23,W_rf_wr_data_22,W_rf_wr_data_21,W_rf_wr_data_20,W_rf_wr_data_19,W_rf_wr_data_18,W_rf_wr_data_17,W_rf_wr_data_16,W_rf_wr_data_15,
W_rf_wr_data_14,W_rf_wr_data_13,W_rf_wr_data_12,W_rf_wr_data_11,W_rf_wr_data_10,W_rf_wr_data_9,W_rf_wr_data_8,W_rf_wr_data_7,W_rf_wr_data_6,W_rf_wr_data_5,W_rf_wr_data_4,W_rf_wr_data_3,W_rf_wr_data_2,W_rf_wr_data_1,W_rf_wr_data_0}),
	.address_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,R_dst_regnum_4,R_dst_regnum_3,R_dst_regnum_2,R_dst_regnum_1,R_dst_regnum_0}),
	.address_b({D_iw_31,D_iw_30,D_iw_29,D_iw_28,D_iw_27}),
	.clock0(clk_clk));

endmodule

module processor_altsyncram_2 (
	q_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[12:0] address_a;
input 	[4:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



processor_altsyncram_vlc1 auto_generated(
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.wren_a(wren_a),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module processor_altsyncram_vlc1 (
	q_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[4:0] address_a;
input 	[4:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

cyclone10lp_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 5;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 31;
defparam ram_block1a4.port_a_logical_ram_depth = 32;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 5;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 31;
defparam ram_block1a4.port_b_logical_ram_depth = 32;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 5;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 31;
defparam ram_block1a3.port_a_logical_ram_depth = 32;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 5;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 31;
defparam ram_block1a3.port_b_logical_ram_depth = 32;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 5;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 31;
defparam ram_block1a2.port_a_logical_ram_depth = 32;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 5;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 31;
defparam ram_block1a2.port_b_logical_ram_depth = 32;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 5;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 31;
defparam ram_block1a1.port_a_logical_ram_depth = 32;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 5;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 31;
defparam ram_block1a1.port_b_logical_ram_depth = 32;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 5;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 31;
defparam ram_block1a0.port_b_logical_ram_depth = 32;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock0";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock0";
defparam ram_block1a16.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus));
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 5;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 31;
defparam ram_block1a31.port_a_logical_ram_depth = 32;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock0";
defparam ram_block1a31.port_b_address_width = 5;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 31;
defparam ram_block1a31.port_b_logical_ram_depth = 32;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock0";
defparam ram_block1a31.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus));
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 5;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 31;
defparam ram_block1a30.port_a_logical_ram_depth = 32;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock0";
defparam ram_block1a30.port_b_address_width = 5;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 31;
defparam ram_block1a30.port_b_logical_ram_depth = 32;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock0";
defparam ram_block1a30.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus));
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 5;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 31;
defparam ram_block1a29.port_a_logical_ram_depth = 32;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock0";
defparam ram_block1a29.port_b_address_width = 5;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 31;
defparam ram_block1a29.port_b_logical_ram_depth = 32;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock0";
defparam ram_block1a29.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus));
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 5;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 31;
defparam ram_block1a28.port_a_logical_ram_depth = 32;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock0";
defparam ram_block1a28.port_b_address_width = 5;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 31;
defparam ram_block1a28.port_b_logical_ram_depth = 32;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock0";
defparam ram_block1a28.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus));
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 5;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 31;
defparam ram_block1a27.port_a_logical_ram_depth = 32;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock0";
defparam ram_block1a27.port_b_address_width = 5;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 31;
defparam ram_block1a27.port_b_logical_ram_depth = 32;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock0";
defparam ram_block1a27.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus));
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 5;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 31;
defparam ram_block1a26.port_a_logical_ram_depth = 32;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock0";
defparam ram_block1a26.port_b_address_width = 5;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 31;
defparam ram_block1a26.port_b_logical_ram_depth = 32;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock0";
defparam ram_block1a26.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus));
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 5;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 31;
defparam ram_block1a25.port_a_logical_ram_depth = 32;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock0";
defparam ram_block1a25.port_b_address_width = 5;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 31;
defparam ram_block1a25.port_b_logical_ram_depth = 32;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock0";
defparam ram_block1a25.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus));
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 5;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 31;
defparam ram_block1a24.port_a_logical_ram_depth = 32;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock0";
defparam ram_block1a24.port_b_address_width = 5;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 31;
defparam ram_block1a24.port_b_logical_ram_depth = 32;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock0";
defparam ram_block1a24.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus));
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 5;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 31;
defparam ram_block1a23.port_a_logical_ram_depth = 32;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock0";
defparam ram_block1a23.port_b_address_width = 5;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 31;
defparam ram_block1a23.port_b_logical_ram_depth = 32;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock0";
defparam ram_block1a23.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus));
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 5;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 31;
defparam ram_block1a22.port_a_logical_ram_depth = 32;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock0";
defparam ram_block1a22.port_b_address_width = 5;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 31;
defparam ram_block1a22.port_b_logical_ram_depth = 32;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock0";
defparam ram_block1a22.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock0";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock0";
defparam ram_block1a21.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock0";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock0";
defparam ram_block1a20.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock0";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock0";
defparam ram_block1a19.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock0";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock0";
defparam ram_block1a18.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_a_module:processor_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock0";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock0";
defparam ram_block1a17.ram_block_type = "auto";

endmodule

module processor_processor_nios2_gen2_0_cpu_register_bank_b_module (
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_16,
	q_b_15,
	q_b_14,
	q_b_13,
	q_b_12,
	q_b_11,
	q_b_10,
	q_b_9,
	q_b_8,
	q_b_31,
	q_b_30,
	q_b_29,
	q_b_28,
	q_b_27,
	q_b_26,
	q_b_25,
	q_b_24,
	q_b_23,
	q_b_22,
	q_b_21,
	q_b_20,
	q_b_19,
	q_b_18,
	q_b_17,
	W_rf_wren,
	W_rf_wr_data_0,
	R_dst_regnum_0,
	R_dst_regnum_1,
	R_dst_regnum_2,
	R_dst_regnum_3,
	R_dst_regnum_4,
	D_iw_22,
	D_iw_23,
	D_iw_24,
	D_iw_25,
	D_iw_26,
	W_rf_wr_data_1,
	W_rf_wr_data_2,
	W_rf_wr_data_3,
	W_rf_wr_data_4,
	W_rf_wr_data_5,
	W_rf_wr_data_6,
	W_rf_wr_data_7,
	W_rf_wr_data_16,
	W_rf_wr_data_15,
	W_rf_wr_data_14,
	W_rf_wr_data_13,
	W_rf_wr_data_12,
	W_rf_wr_data_11,
	W_rf_wr_data_10,
	W_rf_wr_data_9,
	W_rf_wr_data_8,
	W_rf_wr_data_31,
	W_rf_wr_data_30,
	W_rf_wr_data_29,
	W_rf_wr_data_28,
	W_rf_wr_data_27,
	W_rf_wr_data_26,
	W_rf_wr_data_25,
	W_rf_wr_data_24,
	W_rf_wr_data_23,
	W_rf_wr_data_22,
	W_rf_wr_data_21,
	W_rf_wr_data_20,
	W_rf_wr_data_19,
	W_rf_wr_data_18,
	W_rf_wr_data_17,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
output 	q_b_16;
output 	q_b_15;
output 	q_b_14;
output 	q_b_13;
output 	q_b_12;
output 	q_b_11;
output 	q_b_10;
output 	q_b_9;
output 	q_b_8;
output 	q_b_31;
output 	q_b_30;
output 	q_b_29;
output 	q_b_28;
output 	q_b_27;
output 	q_b_26;
output 	q_b_25;
output 	q_b_24;
output 	q_b_23;
output 	q_b_22;
output 	q_b_21;
output 	q_b_20;
output 	q_b_19;
output 	q_b_18;
output 	q_b_17;
input 	W_rf_wren;
input 	W_rf_wr_data_0;
input 	R_dst_regnum_0;
input 	R_dst_regnum_1;
input 	R_dst_regnum_2;
input 	R_dst_regnum_3;
input 	R_dst_regnum_4;
input 	D_iw_22;
input 	D_iw_23;
input 	D_iw_24;
input 	D_iw_25;
input 	D_iw_26;
input 	W_rf_wr_data_1;
input 	W_rf_wr_data_2;
input 	W_rf_wr_data_3;
input 	W_rf_wr_data_4;
input 	W_rf_wr_data_5;
input 	W_rf_wr_data_6;
input 	W_rf_wr_data_7;
input 	W_rf_wr_data_16;
input 	W_rf_wr_data_15;
input 	W_rf_wr_data_14;
input 	W_rf_wr_data_13;
input 	W_rf_wr_data_12;
input 	W_rf_wr_data_11;
input 	W_rf_wr_data_10;
input 	W_rf_wr_data_9;
input 	W_rf_wr_data_8;
input 	W_rf_wr_data_31;
input 	W_rf_wr_data_30;
input 	W_rf_wr_data_29;
input 	W_rf_wr_data_28;
input 	W_rf_wr_data_27;
input 	W_rf_wr_data_26;
input 	W_rf_wr_data_25;
input 	W_rf_wr_data_24;
input 	W_rf_wr_data_23;
input 	W_rf_wr_data_22;
input 	W_rf_wr_data_21;
input 	W_rf_wr_data_20;
input 	W_rf_wr_data_19;
input 	W_rf_wr_data_18;
input 	W_rf_wr_data_17;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



processor_altsyncram_3 the_altsyncram(
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.wren_a(W_rf_wren),
	.data_a({W_rf_wr_data_31,W_rf_wr_data_30,W_rf_wr_data_29,W_rf_wr_data_28,W_rf_wr_data_27,W_rf_wr_data_26,W_rf_wr_data_25,W_rf_wr_data_24,W_rf_wr_data_23,W_rf_wr_data_22,W_rf_wr_data_21,W_rf_wr_data_20,W_rf_wr_data_19,W_rf_wr_data_18,W_rf_wr_data_17,W_rf_wr_data_16,W_rf_wr_data_15,
W_rf_wr_data_14,W_rf_wr_data_13,W_rf_wr_data_12,W_rf_wr_data_11,W_rf_wr_data_10,W_rf_wr_data_9,W_rf_wr_data_8,W_rf_wr_data_7,W_rf_wr_data_6,W_rf_wr_data_5,W_rf_wr_data_4,W_rf_wr_data_3,W_rf_wr_data_2,W_rf_wr_data_1,W_rf_wr_data_0}),
	.address_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,R_dst_regnum_4,R_dst_regnum_3,R_dst_regnum_2,R_dst_regnum_1,R_dst_regnum_0}),
	.address_b({D_iw_26,D_iw_25,D_iw_24,D_iw_23,D_iw_22}),
	.clock0(clk_clk));

endmodule

module processor_altsyncram_3 (
	q_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[12:0] address_a;
input 	[4:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



processor_altsyncram_vlc1_1 auto_generated(
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.wren_a(wren_a),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module processor_altsyncram_vlc1_1 (
	q_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[4:0] address_a;
input 	[4:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

cyclone10lp_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 5;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 31;
defparam ram_block1a0.port_b_logical_ram_depth = 32;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 5;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 31;
defparam ram_block1a1.port_a_logical_ram_depth = 32;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 5;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 31;
defparam ram_block1a1.port_b_logical_ram_depth = 32;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 5;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 31;
defparam ram_block1a2.port_a_logical_ram_depth = 32;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 5;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 31;
defparam ram_block1a2.port_b_logical_ram_depth = 32;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 5;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 31;
defparam ram_block1a3.port_a_logical_ram_depth = 32;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 5;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 31;
defparam ram_block1a3.port_b_logical_ram_depth = 32;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 5;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 31;
defparam ram_block1a4.port_a_logical_ram_depth = 32;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 5;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 31;
defparam ram_block1a4.port_b_logical_ram_depth = 32;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock0";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock0";
defparam ram_block1a16.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus));
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 5;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 31;
defparam ram_block1a31.port_a_logical_ram_depth = 32;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock0";
defparam ram_block1a31.port_b_address_width = 5;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 31;
defparam ram_block1a31.port_b_logical_ram_depth = 32;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock0";
defparam ram_block1a31.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus));
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 5;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 31;
defparam ram_block1a30.port_a_logical_ram_depth = 32;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock0";
defparam ram_block1a30.port_b_address_width = 5;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 31;
defparam ram_block1a30.port_b_logical_ram_depth = 32;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock0";
defparam ram_block1a30.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus));
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 5;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 31;
defparam ram_block1a29.port_a_logical_ram_depth = 32;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock0";
defparam ram_block1a29.port_b_address_width = 5;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 31;
defparam ram_block1a29.port_b_logical_ram_depth = 32;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock0";
defparam ram_block1a29.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus));
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 5;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 31;
defparam ram_block1a28.port_a_logical_ram_depth = 32;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock0";
defparam ram_block1a28.port_b_address_width = 5;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 31;
defparam ram_block1a28.port_b_logical_ram_depth = 32;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock0";
defparam ram_block1a28.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus));
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 5;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 31;
defparam ram_block1a27.port_a_logical_ram_depth = 32;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock0";
defparam ram_block1a27.port_b_address_width = 5;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 31;
defparam ram_block1a27.port_b_logical_ram_depth = 32;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock0";
defparam ram_block1a27.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus));
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 5;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 31;
defparam ram_block1a26.port_a_logical_ram_depth = 32;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock0";
defparam ram_block1a26.port_b_address_width = 5;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 31;
defparam ram_block1a26.port_b_logical_ram_depth = 32;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock0";
defparam ram_block1a26.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus));
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 5;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 31;
defparam ram_block1a25.port_a_logical_ram_depth = 32;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock0";
defparam ram_block1a25.port_b_address_width = 5;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 31;
defparam ram_block1a25.port_b_logical_ram_depth = 32;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock0";
defparam ram_block1a25.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus));
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 5;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 31;
defparam ram_block1a24.port_a_logical_ram_depth = 32;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock0";
defparam ram_block1a24.port_b_address_width = 5;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 31;
defparam ram_block1a24.port_b_logical_ram_depth = 32;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock0";
defparam ram_block1a24.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus));
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 5;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 31;
defparam ram_block1a23.port_a_logical_ram_depth = 32;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock0";
defparam ram_block1a23.port_b_address_width = 5;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 31;
defparam ram_block1a23.port_b_logical_ram_depth = 32;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock0";
defparam ram_block1a23.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus));
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 5;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 31;
defparam ram_block1a22.port_a_logical_ram_depth = 32;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock0";
defparam ram_block1a22.port_b_address_width = 5;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 31;
defparam ram_block1a22.port_b_logical_ram_depth = 32;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock0";
defparam ram_block1a22.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock0";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock0";
defparam ram_block1a21.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock0";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock0";
defparam ram_block1a20.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock0";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock0";
defparam ram_block1a19.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock0";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock0";
defparam ram_block1a18.ram_block_type = "auto";

cyclone10lp_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "processor_nios2_gen2_0:nios2_gen2_0|processor_nios2_gen2_0_cpu:cpu|processor_nios2_gen2_0_cpu_register_bank_b_module:processor_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_vlc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock0";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock0";
defparam ram_block1a17.ram_block_type = "auto";

endmodule

module processor_processor_onchip_memory2_0 (
	q_a_0,
	q_a_22,
	q_a_23,
	q_a_24,
	q_a_25,
	q_a_26,
	q_a_1,
	q_a_4,
	q_a_3,
	q_a_2,
	q_a_5,
	q_a_14,
	q_a_15,
	q_a_11,
	q_a_13,
	q_a_16,
	q_a_12,
	q_a_10,
	q_a_9,
	q_a_8,
	q_a_7,
	q_a_6,
	q_a_21,
	q_a_20,
	q_a_19,
	q_a_18,
	q_a_17,
	q_a_27,
	q_a_28,
	q_a_29,
	q_a_30,
	q_a_31,
	saved_grant_0,
	mem_used_1,
	uav_write,
	WideOr1,
	r_early_rst,
	src_payload,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_46,
	src_data_47,
	src_data_48,
	src_data_49,
	src_data_50,
	src_data_32,
	src_payload1,
	src_data_34,
	src_payload2,
	src_payload3,
	src_data_35,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_data_33,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_22;
output 	q_a_23;
output 	q_a_24;
output 	q_a_25;
output 	q_a_26;
output 	q_a_1;
output 	q_a_4;
output 	q_a_3;
output 	q_a_2;
output 	q_a_5;
output 	q_a_14;
output 	q_a_15;
output 	q_a_11;
output 	q_a_13;
output 	q_a_16;
output 	q_a_12;
output 	q_a_10;
output 	q_a_9;
output 	q_a_8;
output 	q_a_7;
output 	q_a_6;
output 	q_a_21;
output 	q_a_20;
output 	q_a_19;
output 	q_a_18;
output 	q_a_17;
output 	q_a_27;
output 	q_a_28;
output 	q_a_29;
output 	q_a_30;
output 	q_a_31;
input 	saved_grant_0;
input 	mem_used_1;
input 	uav_write;
input 	WideOr1;
input 	r_early_rst;
input 	src_payload;
input 	src_data_38;
input 	src_data_39;
input 	src_data_40;
input 	src_data_41;
input 	src_data_42;
input 	src_data_43;
input 	src_data_44;
input 	src_data_45;
input 	src_data_46;
input 	src_data_47;
input 	src_data_48;
input 	src_data_49;
input 	src_data_50;
input 	src_data_32;
input 	src_payload1;
input 	src_data_34;
input 	src_payload2;
input 	src_payload3;
input 	src_data_35;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_data_33;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wren~0_combout ;


processor_altsyncram_4 the_altsyncram(
	.q_a({q_a_31,q_a_30,q_a_29,q_a_28,q_a_27,q_a_26,q_a_25,q_a_24,q_a_23,q_a_22,q_a_21,q_a_20,q_a_19,q_a_18,q_a_17,q_a_16,q_a_15,q_a_14,q_a_13,q_a_12,q_a_11,q_a_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.clocken0(r_early_rst),
	.wren_a(\wren~0_combout ),
	.data_a({src_payload31,src_payload30,src_payload29,src_payload28,src_payload27,src_payload5,src_payload4,src_payload3,src_payload2,src_payload1,src_payload22,src_payload23,src_payload24,src_payload25,src_payload26,src_payload15,src_payload12,src_payload11,src_payload14,src_payload16,
src_payload13,src_payload17,src_payload18,src_payload19,src_payload20,src_payload21,src_payload10,src_payload7,src_payload8,src_payload9,src_payload6,src_payload}),
	.address_a({src_data_50,src_data_49,src_data_48,src_data_47,src_data_46,src_data_45,src_data_44,src_data_43,src_data_42,src_data_41,src_data_40,src_data_39,src_data_38}),
	.byteena_a({src_data_35,src_data_34,src_data_33,src_data_32}),
	.clock0(clk_clk));

cyclone10lp_lcell_comb \wren~0 (
	.dataa(mem_used_1),
	.datab(uav_write),
	.datac(saved_grant_0),
	.datad(WideOr1),
	.cin(gnd),
	.combout(\wren~0_combout ),
	.cout());
defparam \wren~0 .lut_mask = 16'hBFFF;
defparam \wren~0 .sum_lutc_input = "datac";

endmodule

module processor_altsyncram_4 (
	q_a,
	clocken0,
	wren_a,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	clocken0;
input 	wren_a;
input 	[31:0] data_a;
input 	[12:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



processor_altsyncram_sch1 auto_generated(
	.q_a({q_a[31],q_a[30],q_a[29],q_a[28],q_a[27],q_a[26],q_a[25],q_a[24],q_a[23],q_a[22],q_a[21],q_a[20],q_a[19],q_a[18],q_a[17],q_a[16],q_a[15],q_a[14],q_a[13],q_a[12],q_a[11],q_a[10],q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.clocken0(clocken0),
	.wren_a(wren_a),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.byteena_a({byteena_a[3],byteena_a[2],byteena_a[1],byteena_a[0]}),
	.clock0(clock0));

endmodule

module processor_altsyncram_sch1 (
	q_a,
	clocken0,
	wren_a,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	clocken0;
input 	wren_a;
input 	[31:0] data_a;
input 	[12:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;
wire [143:0] ram_block1a24_PORTADATAOUT_bus;
wire [143:0] ram_block1a25_PORTADATAOUT_bus;
wire [143:0] ram_block1a26_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;
wire [143:0] ram_block1a27_PORTADATAOUT_bus;
wire [143:0] ram_block1a28_PORTADATAOUT_bus;
wire [143:0] ram_block1a29_PORTADATAOUT_bus;
wire [143:0] ram_block1a30_PORTADATAOUT_bus;
wire [143:0] ram_block1a31_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[22] = ram_block1a22_PORTADATAOUT_bus[0];

assign q_a[23] = ram_block1a23_PORTADATAOUT_bus[0];

assign q_a[24] = ram_block1a24_PORTADATAOUT_bus[0];

assign q_a[25] = ram_block1a25_PORTADATAOUT_bus[0];

assign q_a[26] = ram_block1a26_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[14] = ram_block1a14_PORTADATAOUT_bus[0];

assign q_a[15] = ram_block1a15_PORTADATAOUT_bus[0];

assign q_a[11] = ram_block1a11_PORTADATAOUT_bus[0];

assign q_a[13] = ram_block1a13_PORTADATAOUT_bus[0];

assign q_a[16] = ram_block1a16_PORTADATAOUT_bus[0];

assign q_a[12] = ram_block1a12_PORTADATAOUT_bus[0];

assign q_a[10] = ram_block1a10_PORTADATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[21] = ram_block1a21_PORTADATAOUT_bus[0];

assign q_a[20] = ram_block1a20_PORTADATAOUT_bus[0];

assign q_a[19] = ram_block1a19_PORTADATAOUT_bus[0];

assign q_a[18] = ram_block1a18_PORTADATAOUT_bus[0];

assign q_a[17] = ram_block1a17_PORTADATAOUT_bus[0];

assign q_a[27] = ram_block1a27_PORTADATAOUT_bus[0];

assign q_a[28] = ram_block1a28_PORTADATAOUT_bus[0];

assign q_a[29] = ram_block1a29_PORTADATAOUT_bus[0];

assign q_a[30] = ram_block1a30_PORTADATAOUT_bus[0];

assign q_a[31] = ram_block1a31_PORTADATAOUT_bus[0];

cyclone10lp_ram_block ram_block1a0(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "single_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 13;
defparam ram_block1a0.port_a_byte_enable_mask_width = 1;
defparam ram_block1a0.port_a_byte_size = 1;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 8191;
defparam ram_block1a0.port_a_logical_ram_depth = 8192;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a0.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a0.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a0.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a22(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a22.init_file_layout = "port_a";
defparam ram_block1a22.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.operation_mode = "single_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 13;
defparam ram_block1a22.port_a_byte_enable_mask_width = 1;
defparam ram_block1a22.port_a_byte_size = 1;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 8191;
defparam ram_block1a22.port_a_logical_ram_depth = 8192;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.ram_block_type = "auto";
defparam ram_block1a22.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a22.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a22.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a22.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a23(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a23.init_file_layout = "port_a";
defparam ram_block1a23.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.operation_mode = "single_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 13;
defparam ram_block1a23.port_a_byte_enable_mask_width = 1;
defparam ram_block1a23.port_a_byte_size = 1;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 8191;
defparam ram_block1a23.port_a_logical_ram_depth = 8192;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.ram_block_type = "auto";
defparam ram_block1a23.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a23.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a23.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a23.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a24(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a24_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a24.init_file_layout = "port_a";
defparam ram_block1a24.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.operation_mode = "single_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 13;
defparam ram_block1a24.port_a_byte_enable_mask_width = 1;
defparam ram_block1a24.port_a_byte_size = 1;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 8191;
defparam ram_block1a24.port_a_logical_ram_depth = 8192;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.ram_block_type = "auto";
defparam ram_block1a24.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a24.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a24.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a24.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a25(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a25_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a25.init_file_layout = "port_a";
defparam ram_block1a25.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.operation_mode = "single_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 13;
defparam ram_block1a25.port_a_byte_enable_mask_width = 1;
defparam ram_block1a25.port_a_byte_size = 1;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 8191;
defparam ram_block1a25.port_a_logical_ram_depth = 8192;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.ram_block_type = "auto";
defparam ram_block1a25.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a25.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a25.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a25.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a26(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a26_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a26.init_file_layout = "port_a";
defparam ram_block1a26.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.operation_mode = "single_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 13;
defparam ram_block1a26.port_a_byte_enable_mask_width = 1;
defparam ram_block1a26.port_a_byte_size = 1;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 8191;
defparam ram_block1a26.port_a_logical_ram_depth = 8192;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.ram_block_type = "auto";
defparam ram_block1a26.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a26.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a26.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a26.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a1(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "single_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 13;
defparam ram_block1a1.port_a_byte_enable_mask_width = 1;
defparam ram_block1a1.port_a_byte_size = 1;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 8191;
defparam ram_block1a1.port_a_logical_ram_depth = 8192;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a1.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a1.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a1.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a4(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "single_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 13;
defparam ram_block1a4.port_a_byte_enable_mask_width = 1;
defparam ram_block1a4.port_a_byte_size = 1;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 8191;
defparam ram_block1a4.port_a_logical_ram_depth = 8192;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a4.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a4.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a4.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a3(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "single_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 13;
defparam ram_block1a3.port_a_byte_enable_mask_width = 1;
defparam ram_block1a3.port_a_byte_size = 1;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 8191;
defparam ram_block1a3.port_a_logical_ram_depth = 8192;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a3.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a3.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a3.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a2(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "single_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 13;
defparam ram_block1a2.port_a_byte_enable_mask_width = 1;
defparam ram_block1a2.port_a_byte_size = 1;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 8191;
defparam ram_block1a2.port_a_logical_ram_depth = 8192;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a2.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a2.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a2.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a5(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "single_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 13;
defparam ram_block1a5.port_a_byte_enable_mask_width = 1;
defparam ram_block1a5.port_a_byte_size = 1;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 8191;
defparam ram_block1a5.port_a_logical_ram_depth = 8192;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a5.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a5.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a5.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a14(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a14.init_file_layout = "port_a";
defparam ram_block1a14.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.operation_mode = "single_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 13;
defparam ram_block1a14.port_a_byte_enable_mask_width = 1;
defparam ram_block1a14.port_a_byte_size = 1;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 8191;
defparam ram_block1a14.port_a_logical_ram_depth = 8192;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.ram_block_type = "auto";
defparam ram_block1a14.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a14.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a14.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a14.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a15(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a15.init_file_layout = "port_a";
defparam ram_block1a15.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.operation_mode = "single_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 13;
defparam ram_block1a15.port_a_byte_enable_mask_width = 1;
defparam ram_block1a15.port_a_byte_size = 1;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 8191;
defparam ram_block1a15.port_a_logical_ram_depth = 8192;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.ram_block_type = "auto";
defparam ram_block1a15.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a15.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a15.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a15.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a11(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a11.init_file_layout = "port_a";
defparam ram_block1a11.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.operation_mode = "single_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 13;
defparam ram_block1a11.port_a_byte_enable_mask_width = 1;
defparam ram_block1a11.port_a_byte_size = 1;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 8191;
defparam ram_block1a11.port_a_logical_ram_depth = 8192;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a11.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a11.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a11.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a13(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a13.init_file_layout = "port_a";
defparam ram_block1a13.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.operation_mode = "single_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 13;
defparam ram_block1a13.port_a_byte_enable_mask_width = 1;
defparam ram_block1a13.port_a_byte_size = 1;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 8191;
defparam ram_block1a13.port_a_logical_ram_depth = 8192;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a13.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a13.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a13.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a16(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a16.init_file_layout = "port_a";
defparam ram_block1a16.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.operation_mode = "single_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 13;
defparam ram_block1a16.port_a_byte_enable_mask_width = 1;
defparam ram_block1a16.port_a_byte_size = 1;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 8191;
defparam ram_block1a16.port_a_logical_ram_depth = 8192;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.ram_block_type = "auto";
defparam ram_block1a16.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a16.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a16.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a16.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a12(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a12.init_file_layout = "port_a";
defparam ram_block1a12.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.operation_mode = "single_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 13;
defparam ram_block1a12.port_a_byte_enable_mask_width = 1;
defparam ram_block1a12.port_a_byte_size = 1;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 8191;
defparam ram_block1a12.port_a_logical_ram_depth = 8192;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a12.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a12.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a12.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a10(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a10.init_file_layout = "port_a";
defparam ram_block1a10.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.operation_mode = "single_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 13;
defparam ram_block1a10.port_a_byte_enable_mask_width = 1;
defparam ram_block1a10.port_a_byte_size = 1;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 8191;
defparam ram_block1a10.port_a_logical_ram_depth = 8192;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a10.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a10.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a10.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a9(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a9.init_file_layout = "port_a";
defparam ram_block1a9.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "single_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 13;
defparam ram_block1a9.port_a_byte_enable_mask_width = 1;
defparam ram_block1a9.port_a_byte_size = 1;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 8191;
defparam ram_block1a9.port_a_logical_ram_depth = 8192;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a9.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a9.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a9.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a8(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a8.init_file_layout = "port_a";
defparam ram_block1a8.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "single_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 13;
defparam ram_block1a8.port_a_byte_enable_mask_width = 1;
defparam ram_block1a8.port_a_byte_size = 1;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 8191;
defparam ram_block1a8.port_a_logical_ram_depth = 8192;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a8.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a8.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a8.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a7(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "single_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 13;
defparam ram_block1a7.port_a_byte_enable_mask_width = 1;
defparam ram_block1a7.port_a_byte_size = 1;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 8191;
defparam ram_block1a7.port_a_logical_ram_depth = 8192;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a7.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a7.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a7.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a6(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "single_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 13;
defparam ram_block1a6.port_a_byte_enable_mask_width = 1;
defparam ram_block1a6.port_a_byte_size = 1;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 8191;
defparam ram_block1a6.port_a_logical_ram_depth = 8192;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a6.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a6.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a6.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a21(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a21.init_file_layout = "port_a";
defparam ram_block1a21.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.operation_mode = "single_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 13;
defparam ram_block1a21.port_a_byte_enable_mask_width = 1;
defparam ram_block1a21.port_a_byte_size = 1;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 8191;
defparam ram_block1a21.port_a_logical_ram_depth = 8192;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.ram_block_type = "auto";
defparam ram_block1a21.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a21.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a21.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a21.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a20(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a20.init_file_layout = "port_a";
defparam ram_block1a20.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.operation_mode = "single_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 13;
defparam ram_block1a20.port_a_byte_enable_mask_width = 1;
defparam ram_block1a20.port_a_byte_size = 1;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 8191;
defparam ram_block1a20.port_a_logical_ram_depth = 8192;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.ram_block_type = "auto";
defparam ram_block1a20.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a20.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a20.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a20.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a19(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a19.init_file_layout = "port_a";
defparam ram_block1a19.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.operation_mode = "single_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 13;
defparam ram_block1a19.port_a_byte_enable_mask_width = 1;
defparam ram_block1a19.port_a_byte_size = 1;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 8191;
defparam ram_block1a19.port_a_logical_ram_depth = 8192;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.ram_block_type = "auto";
defparam ram_block1a19.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a19.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a19.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a19.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a18(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a18.init_file_layout = "port_a";
defparam ram_block1a18.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.operation_mode = "single_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 13;
defparam ram_block1a18.port_a_byte_enable_mask_width = 1;
defparam ram_block1a18.port_a_byte_size = 1;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 8191;
defparam ram_block1a18.port_a_logical_ram_depth = 8192;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.ram_block_type = "auto";
defparam ram_block1a18.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a18.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a18.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a18.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a17(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a17.init_file_layout = "port_a";
defparam ram_block1a17.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.operation_mode = "single_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 13;
defparam ram_block1a17.port_a_byte_enable_mask_width = 1;
defparam ram_block1a17.port_a_byte_size = 1;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 8191;
defparam ram_block1a17.port_a_logical_ram_depth = 8192;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.ram_block_type = "auto";
defparam ram_block1a17.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a17.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a17.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a17.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a27(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a27_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a27.init_file_layout = "port_a";
defparam ram_block1a27.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.operation_mode = "single_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 13;
defparam ram_block1a27.port_a_byte_enable_mask_width = 1;
defparam ram_block1a27.port_a_byte_size = 1;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 8191;
defparam ram_block1a27.port_a_logical_ram_depth = 8192;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.ram_block_type = "auto";
defparam ram_block1a27.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a27.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a27.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a27.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a28(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a28_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a28.init_file_layout = "port_a";
defparam ram_block1a28.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.operation_mode = "single_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 13;
defparam ram_block1a28.port_a_byte_enable_mask_width = 1;
defparam ram_block1a28.port_a_byte_size = 1;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 8191;
defparam ram_block1a28.port_a_logical_ram_depth = 8192;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.ram_block_type = "auto";
defparam ram_block1a28.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a28.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a28.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a28.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a29(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a29_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a29.init_file_layout = "port_a";
defparam ram_block1a29.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.operation_mode = "single_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 13;
defparam ram_block1a29.port_a_byte_enable_mask_width = 1;
defparam ram_block1a29.port_a_byte_size = 1;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 8191;
defparam ram_block1a29.port_a_logical_ram_depth = 8192;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.ram_block_type = "auto";
defparam ram_block1a29.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a29.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a29.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a29.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a30(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a30_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a30.init_file_layout = "port_a";
defparam ram_block1a30.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.operation_mode = "single_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 13;
defparam ram_block1a30.port_a_byte_enable_mask_width = 1;
defparam ram_block1a30.port_a_byte_size = 1;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 8191;
defparam ram_block1a30.port_a_logical_ram_depth = 8192;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.ram_block_type = "auto";
defparam ram_block1a30.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a30.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a30.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a30.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a31(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a31_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.init_file = "processor_onchip_memory2_0.hex";
defparam ram_block1a31.init_file_layout = "port_a";
defparam ram_block1a31.logical_ram_name = "processor_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_sch1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.operation_mode = "single_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 13;
defparam ram_block1a31.port_a_byte_enable_mask_width = 1;
defparam ram_block1a31.port_a_byte_size = 1;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 8191;
defparam ram_block1a31.port_a_logical_ram_depth = 8192;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.ram_block_type = "auto";
defparam ram_block1a31.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a31.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a31.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a31.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

endmodule

module processor_processor_SEG (
	data_out_0,
	data_out_1,
	data_out_2,
	data_out_3,
	data_out_4,
	data_out_5,
	data_out_6,
	data_out_7,
	writedata,
	reset_n,
	read_mux_out,
	read_mux_out1,
	saved_grant_0,
	src_payload,
	saved_grant_1,
	src_valid,
	src_valid1,
	mem_used_1,
	always0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	readdata_0,
	readdata_1,
	readdata_4,
	readdata_3,
	readdata_2,
	readdata_5,
	readdata_7,
	readdata_6,
	clk)/* synthesis synthesis_greybox=1 */;
output 	data_out_0;
output 	data_out_1;
output 	data_out_2;
output 	data_out_3;
output 	data_out_4;
output 	data_out_5;
output 	data_out_6;
output 	data_out_7;
input 	[31:0] writedata;
input 	reset_n;
input 	read_mux_out;
input 	read_mux_out1;
input 	saved_grant_0;
input 	src_payload;
input 	saved_grant_1;
input 	src_valid;
input 	src_valid1;
input 	mem_used_1;
output 	always0;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
output 	readdata_0;
output 	readdata_1;
output 	readdata_4;
output 	readdata_3;
output 	readdata_2;
output 	readdata_5;
output 	readdata_7;
output 	readdata_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Equal0~0_combout ;
wire \always0~1_combout ;


dffeas \data_out[0] (
	.clk(clk),
	.d(writedata[0]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_0),
	.prn(vcc));
defparam \data_out[0] .is_wysiwyg = "true";
defparam \data_out[0] .power_up = "low";

dffeas \data_out[1] (
	.clk(clk),
	.d(writedata[1]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_1),
	.prn(vcc));
defparam \data_out[1] .is_wysiwyg = "true";
defparam \data_out[1] .power_up = "low";

dffeas \data_out[2] (
	.clk(clk),
	.d(writedata[2]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_2),
	.prn(vcc));
defparam \data_out[2] .is_wysiwyg = "true";
defparam \data_out[2] .power_up = "low";

dffeas \data_out[3] (
	.clk(clk),
	.d(writedata[3]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_3),
	.prn(vcc));
defparam \data_out[3] .is_wysiwyg = "true";
defparam \data_out[3] .power_up = "low";

dffeas \data_out[4] (
	.clk(clk),
	.d(writedata[4]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_4),
	.prn(vcc));
defparam \data_out[4] .is_wysiwyg = "true";
defparam \data_out[4] .power_up = "low";

dffeas \data_out[5] (
	.clk(clk),
	.d(writedata[5]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_5),
	.prn(vcc));
defparam \data_out[5] .is_wysiwyg = "true";
defparam \data_out[5] .power_up = "low";

dffeas \data_out[6] (
	.clk(clk),
	.d(writedata[6]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_6),
	.prn(vcc));
defparam \data_out[6] .is_wysiwyg = "true";
defparam \data_out[6] .power_up = "low";

dffeas \data_out[7] (
	.clk(clk),
	.d(writedata[7]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_7),
	.prn(vcc));
defparam \data_out[7] .is_wysiwyg = "true";
defparam \data_out[7] .power_up = "low";

cyclone10lp_lcell_comb \always0~0 (
	.dataa(src_payload),
	.datab(src_valid),
	.datac(src_valid1),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(always0),
	.cout());
defparam \always0~0 .lut_mask = 16'hFEFF;
defparam \always0~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[0] (
	.dataa(data_out_0),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(readdata_0),
	.cout());
defparam \readdata[0] .lut_mask = 16'hAAFF;
defparam \readdata[0] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[1] (
	.dataa(data_out_1),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(readdata_1),
	.cout());
defparam \readdata[1] .lut_mask = 16'hAAFF;
defparam \readdata[1] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[4] (
	.dataa(data_out_4),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(readdata_4),
	.cout());
defparam \readdata[4] .lut_mask = 16'hAAFF;
defparam \readdata[4] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[3] (
	.dataa(data_out_3),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(readdata_3),
	.cout());
defparam \readdata[3] .lut_mask = 16'hAAFF;
defparam \readdata[3] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[2] (
	.dataa(data_out_2),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(readdata_2),
	.cout());
defparam \readdata[2] .lut_mask = 16'hAAFF;
defparam \readdata[2] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[5] (
	.dataa(data_out_5),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(readdata_5),
	.cout());
defparam \readdata[5] .lut_mask = 16'hAAFF;
defparam \readdata[5] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[7] (
	.dataa(data_out_7),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(readdata_7),
	.cout());
defparam \readdata[7] .lut_mask = 16'hAAFF;
defparam \readdata[7] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[6] (
	.dataa(data_out_6),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(readdata_6),
	.cout());
defparam \readdata[6] .lut_mask = 16'hAAFF;
defparam \readdata[6] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal0~0 (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(read_mux_out1),
	.datad(read_mux_out),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hEFFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \always0~1 (
	.dataa(always0),
	.datab(\Equal0~0_combout ),
	.datac(wait_latency_counter_1),
	.datad(wait_latency_counter_0),
	.cin(gnd),
	.combout(\always0~1_combout ),
	.cout());
defparam \always0~1 .lut_mask = 16'hBFFF;
defparam \always0~1 .sum_lutc_input = "datac";

endmodule

module processor_processor_SEG_EN (
	data_out_0,
	data_out_1,
	data_out_2,
	writedata,
	reset_n,
	read_mux_out,
	read_mux_out1,
	saved_grant_0,
	src_payload,
	saved_grant_1,
	src_valid,
	src_valid1,
	mem_used_1,
	always0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	readdata_0,
	readdata_1,
	readdata_2,
	clk)/* synthesis synthesis_greybox=1 */;
output 	data_out_0;
output 	data_out_1;
output 	data_out_2;
input 	[31:0] writedata;
input 	reset_n;
input 	read_mux_out;
input 	read_mux_out1;
input 	saved_grant_0;
input 	src_payload;
input 	saved_grant_1;
input 	src_valid;
input 	src_valid1;
input 	mem_used_1;
output 	always0;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Equal0~0_combout ;
wire \always0~1_combout ;


dffeas \data_out[0] (
	.clk(clk),
	.d(writedata[0]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_0),
	.prn(vcc));
defparam \data_out[0] .is_wysiwyg = "true";
defparam \data_out[0] .power_up = "low";

dffeas \data_out[1] (
	.clk(clk),
	.d(writedata[1]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_1),
	.prn(vcc));
defparam \data_out[1] .is_wysiwyg = "true";
defparam \data_out[1] .power_up = "low";

dffeas \data_out[2] (
	.clk(clk),
	.d(writedata[2]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_2),
	.prn(vcc));
defparam \data_out[2] .is_wysiwyg = "true";
defparam \data_out[2] .power_up = "low";

cyclone10lp_lcell_comb \always0~0 (
	.dataa(src_payload),
	.datab(src_valid),
	.datac(src_valid1),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(always0),
	.cout());
defparam \always0~0 .lut_mask = 16'hFEFF;
defparam \always0~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[0] (
	.dataa(data_out_0),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(readdata_0),
	.cout());
defparam \readdata[0] .lut_mask = 16'hAAFF;
defparam \readdata[0] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[1] (
	.dataa(data_out_1),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(readdata_1),
	.cout());
defparam \readdata[1] .lut_mask = 16'hAAFF;
defparam \readdata[1] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[2] (
	.dataa(data_out_2),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(readdata_2),
	.cout());
defparam \readdata[2] .lut_mask = 16'hAAFF;
defparam \readdata[2] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal0~0 (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(read_mux_out1),
	.datad(read_mux_out),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hEFFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \always0~1 (
	.dataa(always0),
	.datab(\Equal0~0_combout ),
	.datac(wait_latency_counter_1),
	.datad(wait_latency_counter_0),
	.cin(gnd),
	.combout(\always0~1_combout ),
	.cout());
defparam \always0~1 .lut_mask = 16'hBFFF;
defparam \always0~1 .sum_lutc_input = "datac";

endmodule

module processor_processor_SW (
	W_alu_result_2,
	W_alu_result_3,
	r_sync_rst,
	F_pc_1,
	F_pc_0,
	read_mux_out,
	read_mux_out1,
	saved_grant_0,
	saved_grant_1,
	readdata_0,
	clk_clk,
	sw_export)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_2;
input 	W_alu_result_3;
input 	r_sync_rst;
input 	F_pc_1;
input 	F_pc_0;
output 	read_mux_out;
output 	read_mux_out1;
input 	saved_grant_0;
input 	saved_grant_1;
output 	readdata_0;
input 	clk_clk;
input 	sw_export;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_mux_out~2_combout ;
wire \read_mux_out~3_combout ;


cyclone10lp_lcell_comb \read_mux_out~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(F_pc_1),
	.datad(F_pc_0),
	.cin(gnd),
	.combout(read_mux_out),
	.cout());
defparam \read_mux_out~0 .lut_mask = 16'h0FFF;
defparam \read_mux_out~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \read_mux_out~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(read_mux_out1),
	.cout());
defparam \read_mux_out~1 .lut_mask = 16'h0FFF;
defparam \read_mux_out~1 .sum_lutc_input = "datac";

dffeas \readdata[0] (
	.clk(clk_clk),
	.d(\read_mux_out~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

cyclone10lp_lcell_comb \read_mux_out~2 (
	.dataa(gnd),
	.datab(F_pc_1),
	.datac(F_pc_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(\read_mux_out~2_combout ),
	.cout());
defparam \read_mux_out~2 .lut_mask = 16'h3FFF;
defparam \read_mux_out~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \read_mux_out~3 (
	.dataa(\read_mux_out~2_combout ),
	.datab(sw_export),
	.datac(read_mux_out1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(\read_mux_out~3_combout ),
	.cout());
defparam \read_mux_out~3 .lut_mask = 16'hFEFF;
defparam \read_mux_out~3 .sum_lutc_input = "datac";

endmodule

module processor_processor_uart_0 (
	txd,
	r_sync_rst,
	mem_used_1,
	wait_latency_counter_1,
	src_payload,
	src_data_38,
	src_data_39,
	src_data_40,
	WideOr1,
	av_begintransfer,
	src_data_56,
	rx_rd_strobe_onset,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	readdata_0,
	irq,
	readdata_1,
	readdata_4,
	readdata_3,
	readdata_2,
	readdata_5,
	readdata_9,
	readdata_8,
	readdata_7,
	readdata_6,
	end_begintransfer,
	src_payload9,
	GND_port,
	clk_clk,
	uart_0_rxd)/* synthesis synthesis_greybox=1 */;
output 	txd;
input 	r_sync_rst;
input 	mem_used_1;
input 	wait_latency_counter_1;
input 	src_payload;
input 	src_data_38;
input 	src_data_39;
input 	src_data_40;
input 	WideOr1;
input 	av_begintransfer;
input 	src_data_56;
output 	rx_rd_strobe_onset;
input 	src_payload1;
input 	src_payload2;
input 	src_payload3;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
output 	readdata_0;
output 	irq;
output 	readdata_1;
output 	readdata_4;
output 	readdata_3;
output 	readdata_2;
output 	readdata_5;
output 	readdata_9;
output 	readdata_8;
output 	readdata_7;
output 	readdata_6;
input 	end_begintransfer;
input 	src_payload9;
input 	GND_port;
input 	clk_clk;
input 	uart_0_rxd;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_processor_uart_0_regs|control_reg[9]~q ;
wire \the_processor_uart_0_tx|tx_wr_strobe_onset~0_combout ;
wire \the_processor_uart_0_regs|tx_data[7]~q ;
wire \the_processor_uart_0_regs|tx_data[6]~q ;
wire \the_processor_uart_0_regs|tx_data[5]~q ;
wire \the_processor_uart_0_regs|tx_data[4]~q ;
wire \the_processor_uart_0_regs|tx_data[3]~q ;
wire \the_processor_uart_0_regs|tx_data[2]~q ;
wire \the_processor_uart_0_regs|tx_data[1]~q ;
wire \the_processor_uart_0_regs|tx_data[0]~q ;
wire \the_processor_uart_0_tx|tx_ready~q ;
wire \the_processor_uart_0_tx|tx_wr_strobe_onset~1_combout ;
wire \the_processor_uart_0_rx|rx_data[0]~q ;
wire \the_processor_uart_0_tx|tx_overrun~q ;
wire \the_processor_uart_0_tx|tx_shift_empty~q ;
wire \the_processor_uart_0_rx|break_detect~q ;
wire \the_processor_uart_0_rx|rx_overrun~q ;
wire \the_processor_uart_0_rx|framing_error~q ;
wire \the_processor_uart_0_rx|rx_char_ready~q ;
wire \the_processor_uart_0_rx|rx_data[1]~q ;
wire \the_processor_uart_0_regs|Equal2~0_combout ;
wire \the_processor_uart_0_rx|rx_data[4]~q ;
wire \the_processor_uart_0_rx|rx_data[3]~q ;
wire \the_processor_uart_0_rx|rx_data[2]~q ;
wire \the_processor_uart_0_rx|rx_data[5]~q ;
wire \the_processor_uart_0_rx|rx_data[7]~q ;
wire \the_processor_uart_0_rx|rx_data[6]~q ;
wire \the_processor_uart_0_regs|status_wr_strobe~combout ;


processor_processor_uart_0_regs the_processor_uart_0_regs(
	.reset_n(r_sync_rst),
	.control_reg_9(\the_processor_uart_0_regs|control_reg[9]~q ),
	.writedata({gnd,gnd,gnd,gnd,gnd,gnd,src_payload,src_payload9,src_payload1,src_payload2,src_payload3,src_payload4,src_payload5,src_payload6,src_payload7,src_payload8}),
	.src_data_38(src_data_38),
	.src_data_39(src_data_39),
	.src_data_40(src_data_40),
	.tx_wr_strobe_onset(\the_processor_uart_0_tx|tx_wr_strobe_onset~0_combout ),
	.tx_data_7(\the_processor_uart_0_regs|tx_data[7]~q ),
	.tx_data_6(\the_processor_uart_0_regs|tx_data[6]~q ),
	.tx_data_5(\the_processor_uart_0_regs|tx_data[5]~q ),
	.tx_data_4(\the_processor_uart_0_regs|tx_data[4]~q ),
	.tx_data_3(\the_processor_uart_0_regs|tx_data[3]~q ),
	.tx_data_2(\the_processor_uart_0_regs|tx_data[2]~q ),
	.tx_data_1(\the_processor_uart_0_regs|tx_data[1]~q ),
	.tx_data_0(\the_processor_uart_0_regs|tx_data[0]~q ),
	.tx_ready(\the_processor_uart_0_tx|tx_ready~q ),
	.tx_wr_strobe_onset1(\the_processor_uart_0_tx|tx_wr_strobe_onset~1_combout ),
	.readdata_0(readdata_0),
	.irq1(irq),
	.readdata_1(readdata_1),
	.readdata_4(readdata_4),
	.readdata_3(readdata_3),
	.readdata_2(readdata_2),
	.readdata_5(readdata_5),
	.readdata_9(readdata_9),
	.readdata_8(readdata_8),
	.readdata_7(readdata_7),
	.readdata_6(readdata_6),
	.rx_data_0(\the_processor_uart_0_rx|rx_data[0]~q ),
	.tx_overrun(\the_processor_uart_0_tx|tx_overrun~q ),
	.tx_shift_empty(\the_processor_uart_0_tx|tx_shift_empty~q ),
	.break_detect(\the_processor_uart_0_rx|break_detect~q ),
	.rx_overrun(\the_processor_uart_0_rx|rx_overrun~q ),
	.framing_error(\the_processor_uart_0_rx|framing_error~q ),
	.rx_char_ready(\the_processor_uart_0_rx|rx_char_ready~q ),
	.rx_data_1(\the_processor_uart_0_rx|rx_data[1]~q ),
	.Equal2(\the_processor_uart_0_regs|Equal2~0_combout ),
	.rx_data_4(\the_processor_uart_0_rx|rx_data[4]~q ),
	.rx_data_3(\the_processor_uart_0_rx|rx_data[3]~q ),
	.rx_data_2(\the_processor_uart_0_rx|rx_data[2]~q ),
	.rx_data_5(\the_processor_uart_0_rx|rx_data[5]~q ),
	.rx_data_7(\the_processor_uart_0_rx|rx_data[7]~q ),
	.rx_data_6(\the_processor_uart_0_rx|rx_data[6]~q ),
	.status_wr_strobe1(\the_processor_uart_0_regs|status_wr_strobe~combout ),
	.clk(clk_clk));

processor_processor_uart_0_rx the_processor_uart_0_rx(
	.r_sync_rst(r_sync_rst),
	.mem_used_1(mem_used_1),
	.src_data_38(src_data_38),
	.src_data_39(src_data_39),
	.src_data_40(src_data_40),
	.WideOr1(WideOr1),
	.src_data_56(src_data_56),
	.rx_rd_strobe_onset(rx_rd_strobe_onset),
	.end_begintransfer(end_begintransfer),
	.rx_data_0(\the_processor_uart_0_rx|rx_data[0]~q ),
	.break_detect1(\the_processor_uart_0_rx|break_detect~q ),
	.rx_overrun1(\the_processor_uart_0_rx|rx_overrun~q ),
	.framing_error1(\the_processor_uart_0_rx|framing_error~q ),
	.rx_char_ready1(\the_processor_uart_0_rx|rx_char_ready~q ),
	.rx_data_1(\the_processor_uart_0_rx|rx_data[1]~q ),
	.rx_data_4(\the_processor_uart_0_rx|rx_data[4]~q ),
	.rx_data_3(\the_processor_uart_0_rx|rx_data[3]~q ),
	.rx_data_2(\the_processor_uart_0_rx|rx_data[2]~q ),
	.rx_data_5(\the_processor_uart_0_rx|rx_data[5]~q ),
	.rx_data_7(\the_processor_uart_0_rx|rx_data[7]~q ),
	.rx_data_6(\the_processor_uart_0_rx|rx_data[6]~q ),
	.status_wr_strobe(\the_processor_uart_0_regs|status_wr_strobe~combout ),
	.clk_clk(clk_clk),
	.uart_0_rxd(uart_0_rxd));

processor_processor_uart_0_tx the_processor_uart_0_tx(
	.txd1(txd),
	.reset_n(r_sync_rst),
	.control_reg_9(\the_processor_uart_0_regs|control_reg[9]~q ),
	.mem_used_1(mem_used_1),
	.wait_latency_counter_1(wait_latency_counter_1),
	.src_data_38(src_data_38),
	.src_data_39(src_data_39),
	.src_data_40(src_data_40),
	.WideOr1(WideOr1),
	.av_begintransfer(av_begintransfer),
	.tx_wr_strobe_onset(\the_processor_uart_0_tx|tx_wr_strobe_onset~0_combout ),
	.tx_data_7(\the_processor_uart_0_regs|tx_data[7]~q ),
	.tx_data_6(\the_processor_uart_0_regs|tx_data[6]~q ),
	.tx_data_5(\the_processor_uart_0_regs|tx_data[5]~q ),
	.tx_data_4(\the_processor_uart_0_regs|tx_data[4]~q ),
	.tx_data_3(\the_processor_uart_0_regs|tx_data[3]~q ),
	.tx_data_2(\the_processor_uart_0_regs|tx_data[2]~q ),
	.tx_data_1(\the_processor_uart_0_regs|tx_data[1]~q ),
	.tx_data_0(\the_processor_uart_0_regs|tx_data[0]~q ),
	.tx_ready1(\the_processor_uart_0_tx|tx_ready~q ),
	.tx_wr_strobe_onset1(\the_processor_uart_0_tx|tx_wr_strobe_onset~1_combout ),
	.end_begintransfer(end_begintransfer),
	.tx_overrun1(\the_processor_uart_0_tx|tx_overrun~q ),
	.tx_shift_empty1(\the_processor_uart_0_tx|tx_shift_empty~q ),
	.Equal2(\the_processor_uart_0_regs|Equal2~0_combout ),
	.status_wr_strobe(\the_processor_uart_0_regs|status_wr_strobe~combout ),
	.GND_port(GND_port),
	.clk(clk_clk));

endmodule

module processor_processor_uart_0_regs (
	reset_n,
	control_reg_9,
	writedata,
	src_data_38,
	src_data_39,
	src_data_40,
	tx_wr_strobe_onset,
	tx_data_7,
	tx_data_6,
	tx_data_5,
	tx_data_4,
	tx_data_3,
	tx_data_2,
	tx_data_1,
	tx_data_0,
	tx_ready,
	tx_wr_strobe_onset1,
	readdata_0,
	irq1,
	readdata_1,
	readdata_4,
	readdata_3,
	readdata_2,
	readdata_5,
	readdata_9,
	readdata_8,
	readdata_7,
	readdata_6,
	rx_data_0,
	tx_overrun,
	tx_shift_empty,
	break_detect,
	rx_overrun,
	framing_error,
	rx_char_ready,
	rx_data_1,
	Equal2,
	rx_data_4,
	rx_data_3,
	rx_data_2,
	rx_data_5,
	rx_data_7,
	rx_data_6,
	status_wr_strobe1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	control_reg_9;
input 	[15:0] writedata;
input 	src_data_38;
input 	src_data_39;
input 	src_data_40;
input 	tx_wr_strobe_onset;
output 	tx_data_7;
output 	tx_data_6;
output 	tx_data_5;
output 	tx_data_4;
output 	tx_data_3;
output 	tx_data_2;
output 	tx_data_1;
output 	tx_data_0;
input 	tx_ready;
input 	tx_wr_strobe_onset1;
output 	readdata_0;
output 	irq1;
output 	readdata_1;
output 	readdata_4;
output 	readdata_3;
output 	readdata_2;
output 	readdata_5;
output 	readdata_9;
output 	readdata_8;
output 	readdata_7;
output 	readdata_6;
input 	rx_data_0;
input 	tx_overrun;
input 	tx_shift_empty;
input 	break_detect;
input 	rx_overrun;
input 	framing_error;
input 	rx_char_ready;
input 	rx_data_1;
output 	Equal2;
input 	rx_data_4;
input 	rx_data_3;
input 	rx_data_2;
input 	rx_data_5;
input 	rx_data_7;
input 	rx_data_6;
output 	status_wr_strobe1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \control_wr_strobe~combout ;
wire \control_reg[0]~q ;
wire \selected_read_data[0]~0_combout ;
wire \selected_read_data[0]~1_combout ;
wire \control_reg[4]~q ;
wire \control_reg[5]~q ;
wire \qualified_irq~0_combout ;
wire \control_reg[3]~q ;
wire \control_reg[2]~q ;
wire \qualified_irq~1_combout ;
wire \control_reg[8]~q ;
wire \status_reg[8]~0_combout ;
wire \qualified_irq~2_combout ;
wire \control_reg[7]~q ;
wire \control_reg[1]~q ;
wire \qualified_irq~3_combout ;
wire \control_reg[6]~q ;
wire \qualified_irq~combout ;
wire \selected_read_data~2_combout ;
wire \Equal0~0_combout ;
wire \Equal3~0_combout ;
wire \selected_read_data[1]~3_combout ;
wire \selected_read_data[1]~4_combout ;
wire \selected_read_data~5_combout ;
wire \selected_read_data[4]~6_combout ;
wire \selected_read_data[4]~7_combout ;
wire \selected_read_data~8_combout ;
wire \selected_read_data[3]~9_combout ;
wire \selected_read_data[3]~10_combout ;
wire \selected_read_data~11_combout ;
wire \selected_read_data[2]~12_combout ;
wire \selected_read_data[2]~13_combout ;
wire \selected_read_data~14_combout ;
wire \selected_read_data[5]~15_combout ;
wire \selected_read_data[5]~16_combout ;
wire \selected_read_data~17_combout ;
wire \selected_read_data[8]~combout ;
wire \selected_read_data~18_combout ;
wire \selected_read_data[7]~19_combout ;
wire \selected_read_data[7]~20_combout ;
wire \selected_read_data~21_combout ;
wire \selected_read_data[6]~22_combout ;
wire \selected_read_data[6]~23_combout ;


dffeas \control_reg[9] (
	.clk(clk),
	.d(writedata[9]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\control_wr_strobe~combout ),
	.q(control_reg_9),
	.prn(vcc));
defparam \control_reg[9] .is_wysiwyg = "true";
defparam \control_reg[9] .power_up = "low";

dffeas \tx_data[7] (
	.clk(clk),
	.d(writedata[7]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(tx_wr_strobe_onset1),
	.q(tx_data_7),
	.prn(vcc));
defparam \tx_data[7] .is_wysiwyg = "true";
defparam \tx_data[7] .power_up = "low";

dffeas \tx_data[6] (
	.clk(clk),
	.d(writedata[6]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(tx_wr_strobe_onset1),
	.q(tx_data_6),
	.prn(vcc));
defparam \tx_data[6] .is_wysiwyg = "true";
defparam \tx_data[6] .power_up = "low";

dffeas \tx_data[5] (
	.clk(clk),
	.d(writedata[5]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(tx_wr_strobe_onset1),
	.q(tx_data_5),
	.prn(vcc));
defparam \tx_data[5] .is_wysiwyg = "true";
defparam \tx_data[5] .power_up = "low";

dffeas \tx_data[4] (
	.clk(clk),
	.d(writedata[4]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(tx_wr_strobe_onset1),
	.q(tx_data_4),
	.prn(vcc));
defparam \tx_data[4] .is_wysiwyg = "true";
defparam \tx_data[4] .power_up = "low";

dffeas \tx_data[3] (
	.clk(clk),
	.d(writedata[3]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(tx_wr_strobe_onset1),
	.q(tx_data_3),
	.prn(vcc));
defparam \tx_data[3] .is_wysiwyg = "true";
defparam \tx_data[3] .power_up = "low";

dffeas \tx_data[2] (
	.clk(clk),
	.d(writedata[2]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(tx_wr_strobe_onset1),
	.q(tx_data_2),
	.prn(vcc));
defparam \tx_data[2] .is_wysiwyg = "true";
defparam \tx_data[2] .power_up = "low";

dffeas \tx_data[1] (
	.clk(clk),
	.d(writedata[1]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(tx_wr_strobe_onset1),
	.q(tx_data_1),
	.prn(vcc));
defparam \tx_data[1] .is_wysiwyg = "true";
defparam \tx_data[1] .power_up = "low";

dffeas \tx_data[0] (
	.clk(clk),
	.d(writedata[0]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(tx_wr_strobe_onset1),
	.q(tx_data_0),
	.prn(vcc));
defparam \tx_data[0] .is_wysiwyg = "true";
defparam \tx_data[0] .power_up = "low";

dffeas \readdata[0] (
	.clk(clk),
	.d(\selected_read_data[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas irq(
	.clk(clk),
	.d(\qualified_irq~combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(irq1),
	.prn(vcc));
defparam irq.is_wysiwyg = "true";
defparam irq.power_up = "low";

dffeas \readdata[1] (
	.clk(clk),
	.d(\selected_read_data[1]~4_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[4] (
	.clk(clk),
	.d(\selected_read_data[4]~7_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk),
	.d(\selected_read_data[3]~10_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk),
	.d(\selected_read_data[2]~13_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[5] (
	.clk(clk),
	.d(\selected_read_data[5]~16_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[9] (
	.clk(clk),
	.d(\selected_read_data~17_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_9),
	.prn(vcc));
defparam \readdata[9] .is_wysiwyg = "true";
defparam \readdata[9] .power_up = "low";

dffeas \readdata[8] (
	.clk(clk),
	.d(\selected_read_data[8]~combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_8),
	.prn(vcc));
defparam \readdata[8] .is_wysiwyg = "true";
defparam \readdata[8] .power_up = "low";

dffeas \readdata[7] (
	.clk(clk),
	.d(\selected_read_data[7]~20_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_7),
	.prn(vcc));
defparam \readdata[7] .is_wysiwyg = "true";
defparam \readdata[7] .power_up = "low";

dffeas \readdata[6] (
	.clk(clk),
	.d(\selected_read_data[6]~23_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

cyclone10lp_lcell_comb \Equal2~0 (
	.dataa(src_data_38),
	.datab(gnd),
	.datac(src_data_40),
	.datad(src_data_39),
	.cin(gnd),
	.combout(Equal2),
	.cout());
defparam \Equal2~0 .lut_mask = 16'hAFFF;
defparam \Equal2~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb status_wr_strobe(
	.dataa(src_data_39),
	.datab(src_data_40),
	.datac(src_data_38),
	.datad(tx_wr_strobe_onset),
	.cin(gnd),
	.combout(status_wr_strobe1),
	.cout());
defparam status_wr_strobe.lut_mask = 16'hFFBF;
defparam status_wr_strobe.sum_lutc_input = "datac";

cyclone10lp_lcell_comb control_wr_strobe(
	.dataa(src_data_38),
	.datab(src_data_39),
	.datac(src_data_40),
	.datad(tx_wr_strobe_onset),
	.cin(gnd),
	.combout(\control_wr_strobe~combout ),
	.cout());
defparam control_wr_strobe.lut_mask = 16'hFFEF;
defparam control_wr_strobe.sum_lutc_input = "datac";

dffeas \control_reg[0] (
	.clk(clk),
	.d(writedata[0]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\control_wr_strobe~combout ),
	.q(\control_reg[0]~q ),
	.prn(vcc));
defparam \control_reg[0] .is_wysiwyg = "true";
defparam \control_reg[0] .power_up = "low";

cyclone10lp_lcell_comb \selected_read_data[0]~0 (
	.dataa(tx_data_0),
	.datab(rx_data_0),
	.datac(src_data_38),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\selected_read_data[0]~0_combout ),
	.cout());
defparam \selected_read_data[0]~0 .lut_mask = 16'hEFFE;
defparam \selected_read_data[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \selected_read_data[0]~1 (
	.dataa(\control_reg[0]~q ),
	.datab(src_data_40),
	.datac(src_data_39),
	.datad(\selected_read_data[0]~0_combout ),
	.cin(gnd),
	.combout(\selected_read_data[0]~1_combout ),
	.cout());
defparam \selected_read_data[0]~1 .lut_mask = 16'hFFBF;
defparam \selected_read_data[0]~1 .sum_lutc_input = "datac";

dffeas \control_reg[4] (
	.clk(clk),
	.d(writedata[4]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\control_wr_strobe~combout ),
	.q(\control_reg[4]~q ),
	.prn(vcc));
defparam \control_reg[4] .is_wysiwyg = "true";
defparam \control_reg[4] .power_up = "low";

dffeas \control_reg[5] (
	.clk(clk),
	.d(writedata[5]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\control_wr_strobe~combout ),
	.q(\control_reg[5]~q ),
	.prn(vcc));
defparam \control_reg[5] .is_wysiwyg = "true";
defparam \control_reg[5] .power_up = "low";

cyclone10lp_lcell_comb \qualified_irq~0 (
	.dataa(tx_overrun),
	.datab(\control_reg[4]~q ),
	.datac(\control_reg[5]~q ),
	.datad(tx_shift_empty),
	.cin(gnd),
	.combout(\qualified_irq~0_combout ),
	.cout());
defparam \qualified_irq~0 .lut_mask = 16'hFEFF;
defparam \qualified_irq~0 .sum_lutc_input = "datac";

dffeas \control_reg[3] (
	.clk(clk),
	.d(writedata[3]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\control_wr_strobe~combout ),
	.q(\control_reg[3]~q ),
	.prn(vcc));
defparam \control_reg[3] .is_wysiwyg = "true";
defparam \control_reg[3] .power_up = "low";

dffeas \control_reg[2] (
	.clk(clk),
	.d(writedata[2]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\control_wr_strobe~combout ),
	.q(\control_reg[2]~q ),
	.prn(vcc));
defparam \control_reg[2] .is_wysiwyg = "true";
defparam \control_reg[2] .power_up = "low";

cyclone10lp_lcell_comb \qualified_irq~1 (
	.dataa(break_detect),
	.datab(rx_overrun),
	.datac(\control_reg[3]~q ),
	.datad(\control_reg[2]~q ),
	.cin(gnd),
	.combout(\qualified_irq~1_combout ),
	.cout());
defparam \qualified_irq~1 .lut_mask = 16'hFFFE;
defparam \qualified_irq~1 .sum_lutc_input = "datac";

dffeas \control_reg[8] (
	.clk(clk),
	.d(writedata[8]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\control_wr_strobe~combout ),
	.q(\control_reg[8]~q ),
	.prn(vcc));
defparam \control_reg[8] .is_wysiwyg = "true";
defparam \control_reg[8] .power_up = "low";

cyclone10lp_lcell_comb \status_reg[8]~0 (
	.dataa(tx_overrun),
	.datab(framing_error),
	.datac(break_detect),
	.datad(rx_overrun),
	.cin(gnd),
	.combout(\status_reg[8]~0_combout ),
	.cout());
defparam \status_reg[8]~0 .lut_mask = 16'hFFFE;
defparam \status_reg[8]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \qualified_irq~2 (
	.dataa(\qualified_irq~0_combout ),
	.datab(\qualified_irq~1_combout ),
	.datac(\control_reg[8]~q ),
	.datad(\status_reg[8]~0_combout ),
	.cin(gnd),
	.combout(\qualified_irq~2_combout ),
	.cout());
defparam \qualified_irq~2 .lut_mask = 16'hFFFE;
defparam \qualified_irq~2 .sum_lutc_input = "datac";

dffeas \control_reg[7] (
	.clk(clk),
	.d(writedata[7]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\control_wr_strobe~combout ),
	.q(\control_reg[7]~q ),
	.prn(vcc));
defparam \control_reg[7] .is_wysiwyg = "true";
defparam \control_reg[7] .power_up = "low";

dffeas \control_reg[1] (
	.clk(clk),
	.d(writedata[1]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\control_wr_strobe~combout ),
	.q(\control_reg[1]~q ),
	.prn(vcc));
defparam \control_reg[1] .is_wysiwyg = "true";
defparam \control_reg[1] .power_up = "low";

cyclone10lp_lcell_comb \qualified_irq~3 (
	.dataa(framing_error),
	.datab(rx_char_ready),
	.datac(\control_reg[7]~q ),
	.datad(\control_reg[1]~q ),
	.cin(gnd),
	.combout(\qualified_irq~3_combout ),
	.cout());
defparam \qualified_irq~3 .lut_mask = 16'hFFFE;
defparam \qualified_irq~3 .sum_lutc_input = "datac";

dffeas \control_reg[6] (
	.clk(clk),
	.d(writedata[6]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\control_wr_strobe~combout ),
	.q(\control_reg[6]~q ),
	.prn(vcc));
defparam \control_reg[6] .is_wysiwyg = "true";
defparam \control_reg[6] .power_up = "low";

cyclone10lp_lcell_comb qualified_irq(
	.dataa(\qualified_irq~2_combout ),
	.datab(\qualified_irq~3_combout ),
	.datac(\control_reg[6]~q ),
	.datad(tx_ready),
	.cin(gnd),
	.combout(\qualified_irq~combout ),
	.cout());
defparam qualified_irq.lut_mask = 16'hFEFF;
defparam qualified_irq.sum_lutc_input = "datac";

cyclone10lp_lcell_comb \selected_read_data~2 (
	.dataa(rx_data_1),
	.datab(src_data_40),
	.datac(src_data_38),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\selected_read_data~2_combout ),
	.cout());
defparam \selected_read_data~2 .lut_mask = 16'hBFFF;
defparam \selected_read_data~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal0~0 (
	.dataa(src_data_38),
	.datab(src_data_39),
	.datac(gnd),
	.datad(src_data_40),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hEEFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal3~0 (
	.dataa(src_data_39),
	.datab(gnd),
	.datac(src_data_40),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\Equal3~0_combout ),
	.cout());
defparam \Equal3~0 .lut_mask = 16'hAFFF;
defparam \Equal3~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \selected_read_data[1]~3 (
	.dataa(\Equal0~0_combout ),
	.datab(framing_error),
	.datac(\Equal3~0_combout ),
	.datad(\control_reg[1]~q ),
	.cin(gnd),
	.combout(\selected_read_data[1]~3_combout ),
	.cout());
defparam \selected_read_data[1]~3 .lut_mask = 16'hFFFE;
defparam \selected_read_data[1]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \selected_read_data[1]~4 (
	.dataa(\selected_read_data~2_combout ),
	.datab(\selected_read_data[1]~3_combout ),
	.datac(tx_data_1),
	.datad(Equal2),
	.cin(gnd),
	.combout(\selected_read_data[1]~4_combout ),
	.cout());
defparam \selected_read_data[1]~4 .lut_mask = 16'hFFFE;
defparam \selected_read_data[1]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \selected_read_data~5 (
	.dataa(rx_data_4),
	.datab(src_data_40),
	.datac(src_data_38),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\selected_read_data~5_combout ),
	.cout());
defparam \selected_read_data~5 .lut_mask = 16'hBFFF;
defparam \selected_read_data~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \selected_read_data[4]~6 (
	.dataa(\Equal0~0_combout ),
	.datab(tx_overrun),
	.datac(\Equal3~0_combout ),
	.datad(\control_reg[4]~q ),
	.cin(gnd),
	.combout(\selected_read_data[4]~6_combout ),
	.cout());
defparam \selected_read_data[4]~6 .lut_mask = 16'hFFFE;
defparam \selected_read_data[4]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \selected_read_data[4]~7 (
	.dataa(\selected_read_data~5_combout ),
	.datab(\selected_read_data[4]~6_combout ),
	.datac(tx_data_4),
	.datad(Equal2),
	.cin(gnd),
	.combout(\selected_read_data[4]~7_combout ),
	.cout());
defparam \selected_read_data[4]~7 .lut_mask = 16'hFFFE;
defparam \selected_read_data[4]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \selected_read_data~8 (
	.dataa(rx_data_3),
	.datab(src_data_40),
	.datac(src_data_38),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\selected_read_data~8_combout ),
	.cout());
defparam \selected_read_data~8 .lut_mask = 16'hBFFF;
defparam \selected_read_data~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \selected_read_data[3]~9 (
	.dataa(\Equal0~0_combout ),
	.datab(rx_overrun),
	.datac(\Equal3~0_combout ),
	.datad(\control_reg[3]~q ),
	.cin(gnd),
	.combout(\selected_read_data[3]~9_combout ),
	.cout());
defparam \selected_read_data[3]~9 .lut_mask = 16'hFFFE;
defparam \selected_read_data[3]~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \selected_read_data[3]~10 (
	.dataa(\selected_read_data~8_combout ),
	.datab(\selected_read_data[3]~9_combout ),
	.datac(tx_data_3),
	.datad(Equal2),
	.cin(gnd),
	.combout(\selected_read_data[3]~10_combout ),
	.cout());
defparam \selected_read_data[3]~10 .lut_mask = 16'hFFFE;
defparam \selected_read_data[3]~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \selected_read_data~11 (
	.dataa(rx_data_2),
	.datab(src_data_40),
	.datac(src_data_38),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\selected_read_data~11_combout ),
	.cout());
defparam \selected_read_data~11 .lut_mask = 16'hBFFF;
defparam \selected_read_data~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \selected_read_data[2]~12 (
	.dataa(\Equal0~0_combout ),
	.datab(break_detect),
	.datac(\Equal3~0_combout ),
	.datad(\control_reg[2]~q ),
	.cin(gnd),
	.combout(\selected_read_data[2]~12_combout ),
	.cout());
defparam \selected_read_data[2]~12 .lut_mask = 16'hFFFE;
defparam \selected_read_data[2]~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \selected_read_data[2]~13 (
	.dataa(\selected_read_data~11_combout ),
	.datab(\selected_read_data[2]~12_combout ),
	.datac(tx_data_2),
	.datad(Equal2),
	.cin(gnd),
	.combout(\selected_read_data[2]~13_combout ),
	.cout());
defparam \selected_read_data[2]~13 .lut_mask = 16'hFFFE;
defparam \selected_read_data[2]~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \selected_read_data~14 (
	.dataa(rx_data_5),
	.datab(src_data_40),
	.datac(src_data_38),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\selected_read_data~14_combout ),
	.cout());
defparam \selected_read_data~14 .lut_mask = 16'hBFFF;
defparam \selected_read_data~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \selected_read_data[5]~15 (
	.dataa(\Equal0~0_combout ),
	.datab(\control_reg[5]~q ),
	.datac(\Equal3~0_combout ),
	.datad(tx_shift_empty),
	.cin(gnd),
	.combout(\selected_read_data[5]~15_combout ),
	.cout());
defparam \selected_read_data[5]~15 .lut_mask = 16'hFEFF;
defparam \selected_read_data[5]~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \selected_read_data[5]~16 (
	.dataa(\selected_read_data~14_combout ),
	.datab(\selected_read_data[5]~15_combout ),
	.datac(tx_data_5),
	.datad(Equal2),
	.cin(gnd),
	.combout(\selected_read_data[5]~16_combout ),
	.cout());
defparam \selected_read_data[5]~16 .lut_mask = 16'hFFFE;
defparam \selected_read_data[5]~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \selected_read_data~17 (
	.dataa(control_reg_9),
	.datab(src_data_38),
	.datac(src_data_39),
	.datad(src_data_40),
	.cin(gnd),
	.combout(\selected_read_data~17_combout ),
	.cout());
defparam \selected_read_data~17 .lut_mask = 16'hFEFF;
defparam \selected_read_data~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \selected_read_data[8] (
	.dataa(\Equal0~0_combout ),
	.datab(\status_reg[8]~0_combout ),
	.datac(\Equal3~0_combout ),
	.datad(\control_reg[8]~q ),
	.cin(gnd),
	.combout(\selected_read_data[8]~combout ),
	.cout());
defparam \selected_read_data[8] .lut_mask = 16'hFFFE;
defparam \selected_read_data[8] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \selected_read_data~18 (
	.dataa(rx_data_7),
	.datab(src_data_40),
	.datac(src_data_38),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\selected_read_data~18_combout ),
	.cout());
defparam \selected_read_data~18 .lut_mask = 16'hBFFF;
defparam \selected_read_data~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \selected_read_data[7]~19 (
	.dataa(\Equal0~0_combout ),
	.datab(rx_char_ready),
	.datac(\Equal3~0_combout ),
	.datad(\control_reg[7]~q ),
	.cin(gnd),
	.combout(\selected_read_data[7]~19_combout ),
	.cout());
defparam \selected_read_data[7]~19 .lut_mask = 16'hFFFE;
defparam \selected_read_data[7]~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \selected_read_data[7]~20 (
	.dataa(\selected_read_data~18_combout ),
	.datab(\selected_read_data[7]~19_combout ),
	.datac(tx_data_7),
	.datad(Equal2),
	.cin(gnd),
	.combout(\selected_read_data[7]~20_combout ),
	.cout());
defparam \selected_read_data[7]~20 .lut_mask = 16'hFFFE;
defparam \selected_read_data[7]~20 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \selected_read_data~21 (
	.dataa(rx_data_6),
	.datab(src_data_40),
	.datac(src_data_38),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\selected_read_data~21_combout ),
	.cout());
defparam \selected_read_data~21 .lut_mask = 16'hBFFF;
defparam \selected_read_data~21 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \selected_read_data[6]~22 (
	.dataa(\Equal0~0_combout ),
	.datab(\control_reg[6]~q ),
	.datac(\Equal3~0_combout ),
	.datad(tx_ready),
	.cin(gnd),
	.combout(\selected_read_data[6]~22_combout ),
	.cout());
defparam \selected_read_data[6]~22 .lut_mask = 16'hFEFF;
defparam \selected_read_data[6]~22 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \selected_read_data[6]~23 (
	.dataa(\selected_read_data~21_combout ),
	.datab(\selected_read_data[6]~22_combout ),
	.datac(tx_data_6),
	.datad(Equal2),
	.cin(gnd),
	.combout(\selected_read_data[6]~23_combout ),
	.cout());
defparam \selected_read_data[6]~23 .lut_mask = 16'hFFFE;
defparam \selected_read_data[6]~23 .sum_lutc_input = "datac";

endmodule

module processor_processor_uart_0_rx (
	r_sync_rst,
	mem_used_1,
	src_data_38,
	src_data_39,
	src_data_40,
	WideOr1,
	src_data_56,
	rx_rd_strobe_onset,
	end_begintransfer,
	rx_data_0,
	break_detect1,
	rx_overrun1,
	framing_error1,
	rx_char_ready1,
	rx_data_1,
	rx_data_4,
	rx_data_3,
	rx_data_2,
	rx_data_5,
	rx_data_7,
	rx_data_6,
	status_wr_strobe,
	clk_clk,
	uart_0_rxd)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	mem_used_1;
input 	src_data_38;
input 	src_data_39;
input 	src_data_40;
input 	WideOr1;
input 	src_data_56;
output 	rx_rd_strobe_onset;
input 	end_begintransfer;
output 	rx_data_0;
output 	break_detect1;
output 	rx_overrun1;
output 	framing_error1;
output 	rx_char_ready1;
output 	rx_data_1;
output 	rx_data_4;
output 	rx_data_3;
output 	rx_data_2;
output 	rx_data_5;
output 	rx_data_7;
output 	rx_data_6;
input 	status_wr_strobe;
input 	clk_clk;
input 	uart_0_rxd;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer|dreg[0]~q ;
wire \delayed_unxsync_rxdxx1~q ;
wire \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[0]~1_combout ;
wire \rxd_edge~combout ;
wire \baud_rate_counter~13_combout ;
wire \baud_rate_counter[0]~q ;
wire \Add0~1_cout ;
wire \Add0~2_combout ;
wire \baud_rate_counter~18_combout ;
wire \baud_rate_counter[1]~q ;
wire \Add0~3 ;
wire \Add0~4_combout ;
wire \baud_rate_counter~12_combout ;
wire \baud_rate_counter[2]~q ;
wire \Add0~5 ;
wire \Add0~6_combout ;
wire \Equal0~2_combout ;
wire \baud_rate_counter~17_combout ;
wire \baud_rate_counter[3]~q ;
wire \Add0~7 ;
wire \Add0~8_combout ;
wire \baud_rate_counter~11_combout ;
wire \baud_rate_counter[4]~q ;
wire \Equal0~1_combout ;
wire \always2~0_combout ;
wire \Add0~9 ;
wire \Add0~10_combout ;
wire \baud_rate_counter~16_combout ;
wire \baud_rate_counter[5]~q ;
wire \Add0~11 ;
wire \Add0~12_combout ;
wire \baud_rate_counter~15_combout ;
wire \baud_rate_counter[6]~q ;
wire \Add0~13 ;
wire \Add0~14_combout ;
wire \baud_rate_counter~10_combout ;
wire \baud_rate_counter[7]~q ;
wire \Add0~15 ;
wire \Add0~16_combout ;
wire \baud_rate_counter~14_combout ;
wire \baud_rate_counter[8]~q ;
wire \Equal0~0_combout ;
wire \baud_clk_en~0_combout ;
wire \baud_clk_en~q ;
wire \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[0]~0_combout ;
wire \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[0]~q ;
wire \always4~0_combout ;
wire \do_start_rx~q ;
wire \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[9]~2_combout ;
wire \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[9]~q ;
wire \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[8]~3_combout ;
wire \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[8]~q ;
wire \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[7]~4_combout ;
wire \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[7]~q ;
wire \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[6]~5_combout ;
wire \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[6]~q ;
wire \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[5]~6_combout ;
wire \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[5]~q ;
wire \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[4]~7_combout ;
wire \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[4]~q ;
wire \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[3]~8_combout ;
wire \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[3]~q ;
wire \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[2]~9_combout ;
wire \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[2]~q ;
wire \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[1]~0_combout ;
wire \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[1]~q ;
wire \delayed_unxrx_in_processxx3~q ;
wire \got_new_char~combout ;
wire \WideOr0~0_combout ;
wire \WideOr0~1_combout ;
wire \WideOr0~2_combout ;
wire \break_detect~0_combout ;
wire \rx_overrun~0_combout ;
wire \framing_error~0_combout ;
wire \framing_error~1_combout ;
wire \rx_char_ready~0_combout ;
wire \rx_rd_strobe_onset~1_combout ;
wire \rx_char_ready~1_combout ;


processor_altera_std_synchronizer_5 the_altera_std_synchronizer(
	.reset_n(r_sync_rst),
	.dreg_0(\the_altera_std_synchronizer|dreg[0]~q ),
	.clk(clk_clk),
	.din(uart_0_rxd));

cyclone10lp_lcell_comb \rx_rd_strobe_onset~0 (
	.dataa(WideOr1),
	.datab(gnd),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(rx_rd_strobe_onset),
	.cout());
defparam \rx_rd_strobe_onset~0 .lut_mask = 16'hAAFF;
defparam \rx_rd_strobe_onset~0 .sum_lutc_input = "datac";

dffeas \rx_data[0] (
	.clk(clk_clk),
	.d(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\got_new_char~combout ),
	.q(rx_data_0),
	.prn(vcc));
defparam \rx_data[0] .is_wysiwyg = "true";
defparam \rx_data[0] .power_up = "low";

dffeas break_detect(
	.clk(clk_clk),
	.d(\break_detect~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(break_detect1),
	.prn(vcc));
defparam break_detect.is_wysiwyg = "true";
defparam break_detect.power_up = "low";

dffeas rx_overrun(
	.clk(clk_clk),
	.d(\rx_overrun~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rx_overrun1),
	.prn(vcc));
defparam rx_overrun.is_wysiwyg = "true";
defparam rx_overrun.power_up = "low";

dffeas framing_error(
	.clk(clk_clk),
	.d(\framing_error~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(framing_error1),
	.prn(vcc));
defparam framing_error.is_wysiwyg = "true";
defparam framing_error.power_up = "low";

dffeas rx_char_ready(
	.clk(clk_clk),
	.d(\rx_char_ready~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rx_char_ready1),
	.prn(vcc));
defparam rx_char_ready.is_wysiwyg = "true";
defparam rx_char_ready.power_up = "low";

dffeas \rx_data[1] (
	.clk(clk_clk),
	.d(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\got_new_char~combout ),
	.q(rx_data_1),
	.prn(vcc));
defparam \rx_data[1] .is_wysiwyg = "true";
defparam \rx_data[1] .power_up = "low";

dffeas \rx_data[4] (
	.clk(clk_clk),
	.d(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\got_new_char~combout ),
	.q(rx_data_4),
	.prn(vcc));
defparam \rx_data[4] .is_wysiwyg = "true";
defparam \rx_data[4] .power_up = "low";

dffeas \rx_data[3] (
	.clk(clk_clk),
	.d(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\got_new_char~combout ),
	.q(rx_data_3),
	.prn(vcc));
defparam \rx_data[3] .is_wysiwyg = "true";
defparam \rx_data[3] .power_up = "low";

dffeas \rx_data[2] (
	.clk(clk_clk),
	.d(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\got_new_char~combout ),
	.q(rx_data_2),
	.prn(vcc));
defparam \rx_data[2] .is_wysiwyg = "true";
defparam \rx_data[2] .power_up = "low";

dffeas \rx_data[5] (
	.clk(clk_clk),
	.d(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\got_new_char~combout ),
	.q(rx_data_5),
	.prn(vcc));
defparam \rx_data[5] .is_wysiwyg = "true";
defparam \rx_data[5] .power_up = "low";

dffeas \rx_data[7] (
	.clk(clk_clk),
	.d(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[8]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\got_new_char~combout ),
	.q(rx_data_7),
	.prn(vcc));
defparam \rx_data[7] .is_wysiwyg = "true";
defparam \rx_data[7] .power_up = "low";

dffeas \rx_data[6] (
	.clk(clk_clk),
	.d(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\got_new_char~combout ),
	.q(rx_data_6),
	.prn(vcc));
defparam \rx_data[6] .is_wysiwyg = "true";
defparam \rx_data[6] .power_up = "low";

dffeas delayed_unxsync_rxdxx1(
	.clk(clk_clk),
	.d(\the_altera_std_synchronizer|dreg[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delayed_unxsync_rxdxx1~q ),
	.prn(vcc));
defparam delayed_unxsync_rxdxx1.is_wysiwyg = "true";
defparam delayed_unxsync_rxdxx1.power_up = "low";

cyclone10lp_lcell_comb \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[0]~1 (
	.dataa(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[1]~q ),
	.datab(\do_start_rx~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[0]~1_combout ),
	.cout());
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[0]~1 .lut_mask = 16'hEEEE;
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[0]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb rxd_edge(
	.dataa(gnd),
	.datab(gnd),
	.datac(\the_altera_std_synchronizer|dreg[0]~q ),
	.datad(\delayed_unxsync_rxdxx1~q ),
	.cin(gnd),
	.combout(\rxd_edge~combout ),
	.cout());
defparam rxd_edge.lut_mask = 16'h0FF0;
defparam rxd_edge.sum_lutc_input = "datac";

cyclone10lp_lcell_comb \baud_rate_counter~13 (
	.dataa(\rxd_edge~combout ),
	.datab(\Equal0~0_combout ),
	.datac(\Equal0~1_combout ),
	.datad(\baud_rate_counter[0]~q ),
	.cin(gnd),
	.combout(\baud_rate_counter~13_combout ),
	.cout());
defparam \baud_rate_counter~13 .lut_mask = 16'hBFFF;
defparam \baud_rate_counter~13 .sum_lutc_input = "datac";

dffeas \baud_rate_counter[0] (
	.clk(clk_clk),
	.d(\baud_rate_counter~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_rate_counter[0]~q ),
	.prn(vcc));
defparam \baud_rate_counter[0] .is_wysiwyg = "true";
defparam \baud_rate_counter[0] .power_up = "low";

cyclone10lp_lcell_comb \Add0~1 (
	.dataa(\baud_rate_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\Add0~1_cout ));
defparam \Add0~1 .lut_mask = 16'h00AA;
defparam \Add0~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Add0~2 (
	.dataa(\baud_rate_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1_cout ),
	.combout(\Add0~2_combout ),
	.cout(\Add0~3 ));
defparam \Add0~2 .lut_mask = 16'h5A5F;
defparam \Add0~2 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \baud_rate_counter~18 (
	.dataa(\the_altera_std_synchronizer|dreg[0]~q ),
	.datab(\delayed_unxsync_rxdxx1~q ),
	.datac(\Add0~2_combout ),
	.datad(\always2~0_combout ),
	.cin(gnd),
	.combout(\baud_rate_counter~18_combout ),
	.cout());
defparam \baud_rate_counter~18 .lut_mask = 16'hF9F6;
defparam \baud_rate_counter~18 .sum_lutc_input = "datac";

dffeas \baud_rate_counter[1] (
	.clk(clk_clk),
	.d(\baud_rate_counter~18_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_rate_counter[1]~q ),
	.prn(vcc));
defparam \baud_rate_counter[1] .is_wysiwyg = "true";
defparam \baud_rate_counter[1] .power_up = "low";

cyclone10lp_lcell_comb \Add0~4 (
	.dataa(\baud_rate_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~3 ),
	.combout(\Add0~4_combout ),
	.cout(\Add0~5 ));
defparam \Add0~4 .lut_mask = 16'h5AAF;
defparam \Add0~4 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \baud_rate_counter~12 (
	.dataa(\Add0~4_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\always2~0_combout ),
	.cin(gnd),
	.combout(\baud_rate_counter~12_combout ),
	.cout());
defparam \baud_rate_counter~12 .lut_mask = 16'hAAFF;
defparam \baud_rate_counter~12 .sum_lutc_input = "datac";

dffeas \baud_rate_counter[2] (
	.clk(clk_clk),
	.d(\baud_rate_counter~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_rate_counter[2]~q ),
	.prn(vcc));
defparam \baud_rate_counter[2] .is_wysiwyg = "true";
defparam \baud_rate_counter[2] .power_up = "low";

cyclone10lp_lcell_comb \Add0~6 (
	.dataa(\baud_rate_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~5 ),
	.combout(\Add0~6_combout ),
	.cout(\Add0~7 ));
defparam \Add0~6 .lut_mask = 16'h5A5F;
defparam \Add0~6 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \Equal0~2 (
	.dataa(\Equal0~0_combout ),
	.datab(\Equal0~1_combout ),
	.datac(gnd),
	.datad(\baud_rate_counter[0]~q ),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
defparam \Equal0~2 .lut_mask = 16'hEEFF;
defparam \Equal0~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \baud_rate_counter~17 (
	.dataa(\the_altera_std_synchronizer|dreg[0]~q ),
	.datab(\delayed_unxsync_rxdxx1~q ),
	.datac(\Add0~6_combout ),
	.datad(\Equal0~2_combout ),
	.cin(gnd),
	.combout(\baud_rate_counter~17_combout ),
	.cout());
defparam \baud_rate_counter~17 .lut_mask = 16'hF6FF;
defparam \baud_rate_counter~17 .sum_lutc_input = "datac";

dffeas \baud_rate_counter[3] (
	.clk(clk_clk),
	.d(\baud_rate_counter~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_rate_counter[3]~q ),
	.prn(vcc));
defparam \baud_rate_counter[3] .is_wysiwyg = "true";
defparam \baud_rate_counter[3] .power_up = "low";

cyclone10lp_lcell_comb \Add0~8 (
	.dataa(\baud_rate_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~7 ),
	.combout(\Add0~8_combout ),
	.cout(\Add0~9 ));
defparam \Add0~8 .lut_mask = 16'h5AAF;
defparam \Add0~8 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \baud_rate_counter~11 (
	.dataa(\always2~0_combout ),
	.datab(\Add0~8_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\baud_rate_counter~11_combout ),
	.cout());
defparam \baud_rate_counter~11 .lut_mask = 16'hEEEE;
defparam \baud_rate_counter~11 .sum_lutc_input = "datac";

dffeas \baud_rate_counter[4] (
	.clk(clk_clk),
	.d(\baud_rate_counter~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_rate_counter[4]~q ),
	.prn(vcc));
defparam \baud_rate_counter[4] .is_wysiwyg = "true";
defparam \baud_rate_counter[4] .power_up = "low";

cyclone10lp_lcell_comb \Equal0~1 (
	.dataa(\baud_rate_counter[4]~q ),
	.datab(\baud_rate_counter[3]~q ),
	.datac(\baud_rate_counter[2]~q ),
	.datad(\baud_rate_counter[1]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'h7FFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \always2~0 (
	.dataa(\rxd_edge~combout ),
	.datab(\Equal0~0_combout ),
	.datac(\Equal0~1_combout ),
	.datad(\baud_rate_counter[0]~q ),
	.cin(gnd),
	.combout(\always2~0_combout ),
	.cout());
defparam \always2~0 .lut_mask = 16'hFEFF;
defparam \always2~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Add0~10 (
	.dataa(\baud_rate_counter[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~9 ),
	.combout(\Add0~10_combout ),
	.cout(\Add0~11 ));
defparam \Add0~10 .lut_mask = 16'h5A5F;
defparam \Add0~10 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \baud_rate_counter~16 (
	.dataa(\the_altera_std_synchronizer|dreg[0]~q ),
	.datab(\delayed_unxsync_rxdxx1~q ),
	.datac(\Add0~10_combout ),
	.datad(\always2~0_combout ),
	.cin(gnd),
	.combout(\baud_rate_counter~16_combout ),
	.cout());
defparam \baud_rate_counter~16 .lut_mask = 16'hF9F6;
defparam \baud_rate_counter~16 .sum_lutc_input = "datac";

dffeas \baud_rate_counter[5] (
	.clk(clk_clk),
	.d(\baud_rate_counter~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_rate_counter[5]~q ),
	.prn(vcc));
defparam \baud_rate_counter[5] .is_wysiwyg = "true";
defparam \baud_rate_counter[5] .power_up = "low";

cyclone10lp_lcell_comb \Add0~12 (
	.dataa(\baud_rate_counter[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~11 ),
	.combout(\Add0~12_combout ),
	.cout(\Add0~13 ));
defparam \Add0~12 .lut_mask = 16'h5AAF;
defparam \Add0~12 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \baud_rate_counter~15 (
	.dataa(\the_altera_std_synchronizer|dreg[0]~q ),
	.datab(\delayed_unxsync_rxdxx1~q ),
	.datac(\Add0~12_combout ),
	.datad(\Equal0~2_combout ),
	.cin(gnd),
	.combout(\baud_rate_counter~15_combout ),
	.cout());
defparam \baud_rate_counter~15 .lut_mask = 16'hF6FF;
defparam \baud_rate_counter~15 .sum_lutc_input = "datac";

dffeas \baud_rate_counter[6] (
	.clk(clk_clk),
	.d(\baud_rate_counter~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_rate_counter[6]~q ),
	.prn(vcc));
defparam \baud_rate_counter[6] .is_wysiwyg = "true";
defparam \baud_rate_counter[6] .power_up = "low";

cyclone10lp_lcell_comb \Add0~14 (
	.dataa(\baud_rate_counter[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~13 ),
	.combout(\Add0~14_combout ),
	.cout(\Add0~15 ));
defparam \Add0~14 .lut_mask = 16'h5A5F;
defparam \Add0~14 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \baud_rate_counter~10 (
	.dataa(\always2~0_combout ),
	.datab(\Add0~14_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\baud_rate_counter~10_combout ),
	.cout());
defparam \baud_rate_counter~10 .lut_mask = 16'hEEEE;
defparam \baud_rate_counter~10 .sum_lutc_input = "datac";

dffeas \baud_rate_counter[7] (
	.clk(clk_clk),
	.d(\baud_rate_counter~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_rate_counter[7]~q ),
	.prn(vcc));
defparam \baud_rate_counter[7] .is_wysiwyg = "true";
defparam \baud_rate_counter[7] .power_up = "low";

cyclone10lp_lcell_comb \Add0~16 (
	.dataa(\baud_rate_counter[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add0~15 ),
	.combout(\Add0~16_combout ),
	.cout());
defparam \Add0~16 .lut_mask = 16'h5A5A;
defparam \Add0~16 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \baud_rate_counter~14 (
	.dataa(\the_altera_std_synchronizer|dreg[0]~q ),
	.datab(\delayed_unxsync_rxdxx1~q ),
	.datac(\Add0~16_combout ),
	.datad(\always2~0_combout ),
	.cin(gnd),
	.combout(\baud_rate_counter~14_combout ),
	.cout());
defparam \baud_rate_counter~14 .lut_mask = 16'hF9F6;
defparam \baud_rate_counter~14 .sum_lutc_input = "datac";

dffeas \baud_rate_counter[8] (
	.clk(clk_clk),
	.d(\baud_rate_counter~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_rate_counter[8]~q ),
	.prn(vcc));
defparam \baud_rate_counter[8] .is_wysiwyg = "true";
defparam \baud_rate_counter[8] .power_up = "low";

cyclone10lp_lcell_comb \Equal0~0 (
	.dataa(\baud_rate_counter[8]~q ),
	.datab(\baud_rate_counter[7]~q ),
	.datac(\baud_rate_counter[6]~q ),
	.datad(\baud_rate_counter[5]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'h7FFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \baud_clk_en~0 (
	.dataa(\Equal0~0_combout ),
	.datab(\Equal0~1_combout ),
	.datac(\rxd_edge~combout ),
	.datad(\baud_rate_counter[0]~q ),
	.cin(gnd),
	.combout(\baud_clk_en~0_combout ),
	.cout());
defparam \baud_clk_en~0 .lut_mask = 16'hEFFF;
defparam \baud_clk_en~0 .sum_lutc_input = "datac";

dffeas baud_clk_en(
	.clk(clk_clk),
	.d(\baud_clk_en~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_clk_en~q ),
	.prn(vcc));
defparam baud_clk_en.is_wysiwyg = "true";
defparam baud_clk_en.power_up = "low";

cyclone10lp_lcell_comb \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[0]~0 (
	.dataa(gnd),
	.datab(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[0]~q ),
	.datac(\baud_clk_en~q ),
	.datad(\do_start_rx~q ),
	.cin(gnd),
	.combout(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[0]~0_combout ),
	.cout());
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[0]~0 .lut_mask = 16'hFFFC;
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[0]~0 .sum_lutc_input = "datac";

dffeas \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[0] (
	.clk(clk_clk),
	.d(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[0]~0_combout ),
	.q(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[0]~q ),
	.prn(vcc));
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[0] .is_wysiwyg = "true";
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[0] .power_up = "low";

cyclone10lp_lcell_comb \always4~0 (
	.dataa(\delayed_unxsync_rxdxx1~q ),
	.datab(gnd),
	.datac(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[0]~q ),
	.datad(\the_altera_std_synchronizer|dreg[0]~q ),
	.cin(gnd),
	.combout(\always4~0_combout ),
	.cout());
defparam \always4~0 .lut_mask = 16'hAFFF;
defparam \always4~0 .sum_lutc_input = "datac";

dffeas do_start_rx(
	.clk(clk_clk),
	.d(\always4~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\do_start_rx~q ),
	.prn(vcc));
defparam do_start_rx.is_wysiwyg = "true";
defparam do_start_rx.power_up = "low";

cyclone10lp_lcell_comb \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[9]~2 (
	.dataa(\do_start_rx~q ),
	.datab(\the_altera_std_synchronizer|dreg[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[9]~2_combout ),
	.cout());
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[9]~2 .lut_mask = 16'hEEEE;
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[9]~2 .sum_lutc_input = "datac";

dffeas \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[9] (
	.clk(clk_clk),
	.d(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[9]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[0]~0_combout ),
	.q(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[9]~q ),
	.prn(vcc));
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[9] .is_wysiwyg = "true";
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[9] .power_up = "low";

cyclone10lp_lcell_comb \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[8]~3 (
	.dataa(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[9]~q ),
	.datab(\do_start_rx~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[8]~3_combout ),
	.cout());
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[8]~3 .lut_mask = 16'hEEEE;
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[8]~3 .sum_lutc_input = "datac";

dffeas \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[8] (
	.clk(clk_clk),
	.d(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[8]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[0]~0_combout ),
	.q(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[8]~q ),
	.prn(vcc));
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[8] .is_wysiwyg = "true";
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[8] .power_up = "low";

cyclone10lp_lcell_comb \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[7]~4 (
	.dataa(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[8]~q ),
	.datab(\do_start_rx~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[7]~4_combout ),
	.cout());
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[7]~4 .lut_mask = 16'hEEEE;
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[7]~4 .sum_lutc_input = "datac";

dffeas \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[7] (
	.clk(clk_clk),
	.d(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[7]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[0]~0_combout ),
	.q(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[7]~q ),
	.prn(vcc));
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[7] .is_wysiwyg = "true";
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[7] .power_up = "low";

cyclone10lp_lcell_comb \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[6]~5 (
	.dataa(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[7]~q ),
	.datab(\do_start_rx~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[6]~5_combout ),
	.cout());
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[6]~5 .lut_mask = 16'hEEEE;
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[6]~5 .sum_lutc_input = "datac";

dffeas \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[6] (
	.clk(clk_clk),
	.d(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[6]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[0]~0_combout ),
	.q(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[6]~q ),
	.prn(vcc));
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[6] .is_wysiwyg = "true";
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[6] .power_up = "low";

cyclone10lp_lcell_comb \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[5]~6 (
	.dataa(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[6]~q ),
	.datab(\do_start_rx~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[5]~6_combout ),
	.cout());
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[5]~6 .lut_mask = 16'hEEEE;
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[5]~6 .sum_lutc_input = "datac";

dffeas \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[5] (
	.clk(clk_clk),
	.d(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[5]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[0]~0_combout ),
	.q(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[5]~q ),
	.prn(vcc));
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[5] .is_wysiwyg = "true";
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[5] .power_up = "low";

cyclone10lp_lcell_comb \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[4]~7 (
	.dataa(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[5]~q ),
	.datab(\do_start_rx~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[4]~7_combout ),
	.cout());
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[4]~7 .lut_mask = 16'hEEEE;
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[4]~7 .sum_lutc_input = "datac";

dffeas \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[4] (
	.clk(clk_clk),
	.d(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[4]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[0]~0_combout ),
	.q(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[4]~q ),
	.prn(vcc));
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[4] .is_wysiwyg = "true";
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[4] .power_up = "low";

cyclone10lp_lcell_comb \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[3]~8 (
	.dataa(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[4]~q ),
	.datab(\do_start_rx~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[3]~8_combout ),
	.cout());
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[3]~8 .lut_mask = 16'hEEEE;
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[3]~8 .sum_lutc_input = "datac";

dffeas \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[3] (
	.clk(clk_clk),
	.d(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[3]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[0]~0_combout ),
	.q(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[3]~q ),
	.prn(vcc));
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[3] .is_wysiwyg = "true";
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[3] .power_up = "low";

cyclone10lp_lcell_comb \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[2]~9 (
	.dataa(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[3]~q ),
	.datab(\do_start_rx~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[2]~9_combout ),
	.cout());
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[2]~9 .lut_mask = 16'hEEEE;
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[2]~9 .sum_lutc_input = "datac";

dffeas \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[2] (
	.clk(clk_clk),
	.d(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[2]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[0]~0_combout ),
	.q(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[2]~q ),
	.prn(vcc));
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[2] .is_wysiwyg = "true";
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[2] .power_up = "low";

cyclone10lp_lcell_comb \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[1]~0 (
	.dataa(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[2]~q ),
	.datab(\do_start_rx~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[1]~0_combout ),
	.cout());
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[1]~0 .lut_mask = 16'hEEEE;
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[1]~0 .sum_lutc_input = "datac";

dffeas \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[1] (
	.clk(clk_clk),
	.d(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_in[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[0]~0_combout ),
	.q(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[1]~q ),
	.prn(vcc));
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[1] .is_wysiwyg = "true";
defparam \unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[1] .power_up = "low";

dffeas delayed_unxrx_in_processxx3(
	.clk(clk_clk),
	.d(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delayed_unxrx_in_processxx3~q ),
	.prn(vcc));
defparam delayed_unxrx_in_processxx3.is_wysiwyg = "true";
defparam delayed_unxrx_in_processxx3.power_up = "low";

cyclone10lp_lcell_comb got_new_char(
	.dataa(\delayed_unxrx_in_processxx3~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[0]~q ),
	.cin(gnd),
	.combout(\got_new_char~combout ),
	.cout());
defparam got_new_char.lut_mask = 16'hAAFF;
defparam got_new_char.sum_lutc_input = "datac";

cyclone10lp_lcell_comb \WideOr0~0 (
	.dataa(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[0]~q ),
	.datab(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[9]~q ),
	.datac(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[8]~q ),
	.datad(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[7]~q ),
	.cin(gnd),
	.combout(\WideOr0~0_combout ),
	.cout());
defparam \WideOr0~0 .lut_mask = 16'hFFFE;
defparam \WideOr0~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \WideOr0~1 (
	.dataa(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[6]~q ),
	.datab(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[5]~q ),
	.datac(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[4]~q ),
	.datad(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[3]~q ),
	.cin(gnd),
	.combout(\WideOr0~1_combout ),
	.cout());
defparam \WideOr0~1 .lut_mask = 16'hFFFE;
defparam \WideOr0~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \WideOr0~2 (
	.dataa(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[1]~q ),
	.datab(\WideOr0~0_combout ),
	.datac(\WideOr0~1_combout ),
	.datad(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[2]~q ),
	.cin(gnd),
	.combout(\WideOr0~2_combout ),
	.cout());
defparam \WideOr0~2 .lut_mask = 16'hFFFE;
defparam \WideOr0~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \break_detect~0 (
	.dataa(break_detect1),
	.datab(\got_new_char~combout ),
	.datac(\WideOr0~2_combout ),
	.datad(status_wr_strobe),
	.cin(gnd),
	.combout(\break_detect~0_combout ),
	.cout());
defparam \break_detect~0 .lut_mask = 16'hEFFF;
defparam \break_detect~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \rx_overrun~0 (
	.dataa(rx_overrun1),
	.datab(rx_char_ready1),
	.datac(\got_new_char~combout ),
	.datad(status_wr_strobe),
	.cin(gnd),
	.combout(\rx_overrun~0_combout ),
	.cout());
defparam \rx_overrun~0 .lut_mask = 16'hFEFF;
defparam \rx_overrun~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \framing_error~0 (
	.dataa(\delayed_unxrx_in_processxx3~q ),
	.datab(gnd),
	.datac(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[0]~q ),
	.datad(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[9]~q ),
	.cin(gnd),
	.combout(\framing_error~0_combout ),
	.cout());
defparam \framing_error~0 .lut_mask = 16'hAFFF;
defparam \framing_error~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \framing_error~1 (
	.dataa(framing_error1),
	.datab(\WideOr0~2_combout ),
	.datac(\framing_error~0_combout ),
	.datad(status_wr_strobe),
	.cin(gnd),
	.combout(\framing_error~1_combout ),
	.cout());
defparam \framing_error~1 .lut_mask = 16'hFEFF;
defparam \framing_error~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \rx_char_ready~0 (
	.dataa(rx_char_ready1),
	.datab(\delayed_unxrx_in_processxx3~q ),
	.datac(gnd),
	.datad(\unxshiftxrxd_shift_regxshift_reg_start_bit_nxx6_out[0]~q ),
	.cin(gnd),
	.combout(\rx_char_ready~0_combout ),
	.cout());
defparam \rx_char_ready~0 .lut_mask = 16'hEEFF;
defparam \rx_char_ready~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \rx_rd_strobe_onset~1 (
	.dataa(src_data_40),
	.datab(src_data_38),
	.datac(src_data_39),
	.datad(end_begintransfer),
	.cin(gnd),
	.combout(\rx_rd_strobe_onset~1_combout ),
	.cout());
defparam \rx_rd_strobe_onset~1 .lut_mask = 16'h7FFF;
defparam \rx_rd_strobe_onset~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \rx_char_ready~1 (
	.dataa(\rx_char_ready~0_combout ),
	.datab(rx_rd_strobe_onset),
	.datac(src_data_56),
	.datad(\rx_rd_strobe_onset~1_combout ),
	.cin(gnd),
	.combout(\rx_char_ready~1_combout ),
	.cout());
defparam \rx_char_ready~1 .lut_mask = 16'hBFFF;
defparam \rx_char_ready~1 .sum_lutc_input = "datac";

endmodule

module processor_altera_std_synchronizer_5 (
	reset_n,
	dreg_0,
	clk,
	din)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_0;
input 	clk;
input 	din;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module processor_processor_uart_0_tx (
	txd1,
	reset_n,
	control_reg_9,
	mem_used_1,
	wait_latency_counter_1,
	src_data_38,
	src_data_39,
	src_data_40,
	WideOr1,
	av_begintransfer,
	tx_wr_strobe_onset,
	tx_data_7,
	tx_data_6,
	tx_data_5,
	tx_data_4,
	tx_data_3,
	tx_data_2,
	tx_data_1,
	tx_data_0,
	tx_ready1,
	tx_wr_strobe_onset1,
	end_begintransfer,
	tx_overrun1,
	tx_shift_empty1,
	Equal2,
	status_wr_strobe,
	GND_port,
	clk)/* synthesis synthesis_greybox=1 */;
output 	txd1;
input 	reset_n;
input 	control_reg_9;
input 	mem_used_1;
input 	wait_latency_counter_1;
input 	src_data_38;
input 	src_data_39;
input 	src_data_40;
input 	WideOr1;
input 	av_begintransfer;
output 	tx_wr_strobe_onset;
input 	tx_data_7;
input 	tx_data_6;
input 	tx_data_5;
input 	tx_data_4;
input 	tx_data_3;
input 	tx_data_2;
input 	tx_data_1;
input 	tx_data_0;
output 	tx_ready1;
output 	tx_wr_strobe_onset1;
input 	end_begintransfer;
output 	tx_overrun1;
output 	tx_shift_empty1;
input 	Equal2;
input 	status_wr_strobe;
input 	GND_port;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \pre_txd~0_combout ;
wire \pre_txd~1_combout ;
wire \WideOr0~combout ;
wire \do_load_shifter~0_combout ;
wire \do_load_shifter~q ;
wire \baud_rate_counter[0]~9_combout ;
wire \baud_rate_counter[0]~10 ;
wire \baud_rate_counter[1]~11_combout ;
wire \baud_rate_counter[1]~q ;
wire \baud_rate_counter[1]~12 ;
wire \baud_rate_counter[2]~13_combout ;
wire \baud_rate_counter[2]~q ;
wire \baud_rate_counter[2]~14 ;
wire \baud_rate_counter[3]~15_combout ;
wire \baud_rate_counter[3]~q ;
wire \baud_rate_counter[3]~16 ;
wire \baud_rate_counter[4]~17_combout ;
wire \baud_rate_counter[4]~q ;
wire \baud_rate_counter[4]~18 ;
wire \baud_rate_counter[5]~19_combout ;
wire \baud_rate_counter[5]~q ;
wire \baud_rate_counter[5]~20 ;
wire \baud_rate_counter[6]~21_combout ;
wire \baud_rate_counter[6]~q ;
wire \baud_rate_counter[6]~22 ;
wire \baud_rate_counter[7]~23_combout ;
wire \baud_rate_counter[7]~q ;
wire \Equal0~1_combout ;
wire \baud_rate_counter[7]~24 ;
wire \baud_rate_counter[8]~25_combout ;
wire \baud_rate_counter[8]~q ;
wire \always4~0_combout ;
wire \baud_rate_counter[0]~q ;
wire \Equal0~0_combout ;
wire \Equal0~2_combout ;
wire \baud_clk_en~q ;
wire \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[9]~3_combout ;
wire \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[9]~q ;
wire \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[8]~4_combout ;
wire \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[4]~1_combout ;
wire \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[8]~q ;
wire \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[7]~5_combout ;
wire \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[7]~q ;
wire \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[6]~6_combout ;
wire \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[6]~q ;
wire \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[5]~7_combout ;
wire \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[5]~q ;
wire \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[4]~8_combout ;
wire \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[4]~q ;
wire \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[3]~9_combout ;
wire \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[3]~q ;
wire \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[2]~10_combout ;
wire \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[2]~q ;
wire \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[1]~11_combout ;
wire \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[1]~q ;
wire \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[0]~0_combout ;
wire \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[0]~2_combout ;
wire \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[0]~q ;
wire \pre_txd~2_combout ;
wire \pre_txd~3_combout ;
wire \pre_txd~q ;
wire \txd~0_combout ;
wire \tx_ready~0_combout ;
wire \tx_overrun~0_combout ;
wire \tx_overrun~1_combout ;
wire \tx_shift_empty~0_combout ;


dffeas txd(
	.clk(clk),
	.d(\txd~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(txd1),
	.prn(vcc));
defparam txd.is_wysiwyg = "true";
defparam txd.power_up = "low";

cyclone10lp_lcell_comb \tx_wr_strobe_onset~0 (
	.dataa(WideOr1),
	.datab(av_begintransfer),
	.datac(mem_used_1),
	.datad(wait_latency_counter_1),
	.cin(gnd),
	.combout(tx_wr_strobe_onset),
	.cout());
defparam \tx_wr_strobe_onset~0 .lut_mask = 16'hEFFF;
defparam \tx_wr_strobe_onset~0 .sum_lutc_input = "datac";

dffeas tx_ready(
	.clk(clk),
	.d(\tx_ready~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(tx_ready1),
	.prn(vcc));
defparam tx_ready.is_wysiwyg = "true";
defparam tx_ready.power_up = "low";

cyclone10lp_lcell_comb \tx_wr_strobe_onset~1 (
	.dataa(src_data_38),
	.datab(tx_wr_strobe_onset),
	.datac(src_data_40),
	.datad(src_data_39),
	.cin(gnd),
	.combout(tx_wr_strobe_onset1),
	.cout());
defparam \tx_wr_strobe_onset~1 .lut_mask = 16'hEFFF;
defparam \tx_wr_strobe_onset~1 .sum_lutc_input = "datac";

dffeas tx_overrun(
	.clk(clk),
	.d(\tx_overrun~1_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(tx_overrun1),
	.prn(vcc));
defparam tx_overrun.is_wysiwyg = "true";
defparam tx_overrun.power_up = "low";

dffeas tx_shift_empty(
	.clk(clk),
	.d(\tx_shift_empty~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(tx_shift_empty1),
	.prn(vcc));
defparam tx_shift_empty.is_wysiwyg = "true";
defparam tx_shift_empty.power_up = "low";

cyclone10lp_lcell_comb \pre_txd~0 (
	.dataa(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[9]~q ),
	.datab(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[8]~q ),
	.datac(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[7]~q ),
	.datad(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[6]~q ),
	.cin(gnd),
	.combout(\pre_txd~0_combout ),
	.cout());
defparam \pre_txd~0 .lut_mask = 16'h7FFF;
defparam \pre_txd~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_txd~1 (
	.dataa(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[5]~q ),
	.datab(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[4]~q ),
	.datac(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[3]~q ),
	.datad(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[2]~q ),
	.cin(gnd),
	.combout(\pre_txd~1_combout ),
	.cout());
defparam \pre_txd~1 .lut_mask = 16'h7FFF;
defparam \pre_txd~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb WideOr0(
	.dataa(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[0]~q ),
	.datab(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[1]~q ),
	.datac(\pre_txd~0_combout ),
	.datad(\pre_txd~1_combout ),
	.cin(gnd),
	.combout(\WideOr0~combout ),
	.cout());
defparam WideOr0.lut_mask = 16'hEFFF;
defparam WideOr0.sum_lutc_input = "datac";

cyclone10lp_lcell_comb \do_load_shifter~0 (
	.dataa(\WideOr0~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(tx_ready1),
	.cin(gnd),
	.combout(\do_load_shifter~0_combout ),
	.cout());
defparam \do_load_shifter~0 .lut_mask = 16'hFF55;
defparam \do_load_shifter~0 .sum_lutc_input = "datac";

dffeas do_load_shifter(
	.clk(clk),
	.d(\do_load_shifter~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\do_load_shifter~q ),
	.prn(vcc));
defparam do_load_shifter.is_wysiwyg = "true";
defparam do_load_shifter.power_up = "low";

cyclone10lp_lcell_comb \baud_rate_counter[0]~9 (
	.dataa(\baud_rate_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\baud_rate_counter[0]~9_combout ),
	.cout(\baud_rate_counter[0]~10 ));
defparam \baud_rate_counter[0]~9 .lut_mask = 16'h55AA;
defparam \baud_rate_counter[0]~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \baud_rate_counter[1]~11 (
	.dataa(\baud_rate_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_rate_counter[0]~10 ),
	.combout(\baud_rate_counter[1]~11_combout ),
	.cout(\baud_rate_counter[1]~12 ));
defparam \baud_rate_counter[1]~11 .lut_mask = 16'h5A5F;
defparam \baud_rate_counter[1]~11 .sum_lutc_input = "cin";

dffeas \baud_rate_counter[1] (
	.clk(clk),
	.d(\baud_rate_counter[1]~11_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always4~0_combout ),
	.ena(vcc),
	.q(\baud_rate_counter[1]~q ),
	.prn(vcc));
defparam \baud_rate_counter[1] .is_wysiwyg = "true";
defparam \baud_rate_counter[1] .power_up = "low";

cyclone10lp_lcell_comb \baud_rate_counter[2]~13 (
	.dataa(\baud_rate_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_rate_counter[1]~12 ),
	.combout(\baud_rate_counter[2]~13_combout ),
	.cout(\baud_rate_counter[2]~14 ));
defparam \baud_rate_counter[2]~13 .lut_mask = 16'h5AAF;
defparam \baud_rate_counter[2]~13 .sum_lutc_input = "cin";

dffeas \baud_rate_counter[2] (
	.clk(clk),
	.d(\baud_rate_counter[2]~13_combout ),
	.asdata(GND_port),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always4~0_combout ),
	.ena(vcc),
	.q(\baud_rate_counter[2]~q ),
	.prn(vcc));
defparam \baud_rate_counter[2] .is_wysiwyg = "true";
defparam \baud_rate_counter[2] .power_up = "low";

cyclone10lp_lcell_comb \baud_rate_counter[3]~15 (
	.dataa(\baud_rate_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_rate_counter[2]~14 ),
	.combout(\baud_rate_counter[3]~15_combout ),
	.cout(\baud_rate_counter[3]~16 ));
defparam \baud_rate_counter[3]~15 .lut_mask = 16'h5A5F;
defparam \baud_rate_counter[3]~15 .sum_lutc_input = "cin";

dffeas \baud_rate_counter[3] (
	.clk(clk),
	.d(\baud_rate_counter[3]~15_combout ),
	.asdata(GND_port),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always4~0_combout ),
	.ena(vcc),
	.q(\baud_rate_counter[3]~q ),
	.prn(vcc));
defparam \baud_rate_counter[3] .is_wysiwyg = "true";
defparam \baud_rate_counter[3] .power_up = "low";

cyclone10lp_lcell_comb \baud_rate_counter[4]~17 (
	.dataa(\baud_rate_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_rate_counter[3]~16 ),
	.combout(\baud_rate_counter[4]~17_combout ),
	.cout(\baud_rate_counter[4]~18 ));
defparam \baud_rate_counter[4]~17 .lut_mask = 16'h5AAF;
defparam \baud_rate_counter[4]~17 .sum_lutc_input = "cin";

dffeas \baud_rate_counter[4] (
	.clk(clk),
	.d(\baud_rate_counter[4]~17_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always4~0_combout ),
	.ena(vcc),
	.q(\baud_rate_counter[4]~q ),
	.prn(vcc));
defparam \baud_rate_counter[4] .is_wysiwyg = "true";
defparam \baud_rate_counter[4] .power_up = "low";

cyclone10lp_lcell_comb \baud_rate_counter[5]~19 (
	.dataa(\baud_rate_counter[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_rate_counter[4]~18 ),
	.combout(\baud_rate_counter[5]~19_combout ),
	.cout(\baud_rate_counter[5]~20 ));
defparam \baud_rate_counter[5]~19 .lut_mask = 16'h5A5F;
defparam \baud_rate_counter[5]~19 .sum_lutc_input = "cin";

dffeas \baud_rate_counter[5] (
	.clk(clk),
	.d(\baud_rate_counter[5]~19_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always4~0_combout ),
	.ena(vcc),
	.q(\baud_rate_counter[5]~q ),
	.prn(vcc));
defparam \baud_rate_counter[5] .is_wysiwyg = "true";
defparam \baud_rate_counter[5] .power_up = "low";

cyclone10lp_lcell_comb \baud_rate_counter[6]~21 (
	.dataa(\baud_rate_counter[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_rate_counter[5]~20 ),
	.combout(\baud_rate_counter[6]~21_combout ),
	.cout(\baud_rate_counter[6]~22 ));
defparam \baud_rate_counter[6]~21 .lut_mask = 16'h5AAF;
defparam \baud_rate_counter[6]~21 .sum_lutc_input = "cin";

dffeas \baud_rate_counter[6] (
	.clk(clk),
	.d(\baud_rate_counter[6]~21_combout ),
	.asdata(GND_port),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always4~0_combout ),
	.ena(vcc),
	.q(\baud_rate_counter[6]~q ),
	.prn(vcc));
defparam \baud_rate_counter[6] .is_wysiwyg = "true";
defparam \baud_rate_counter[6] .power_up = "low";

cyclone10lp_lcell_comb \baud_rate_counter[7]~23 (
	.dataa(\baud_rate_counter[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_rate_counter[6]~22 ),
	.combout(\baud_rate_counter[7]~23_combout ),
	.cout(\baud_rate_counter[7]~24 ));
defparam \baud_rate_counter[7]~23 .lut_mask = 16'h5A5F;
defparam \baud_rate_counter[7]~23 .sum_lutc_input = "cin";

dffeas \baud_rate_counter[7] (
	.clk(clk),
	.d(\baud_rate_counter[7]~23_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always4~0_combout ),
	.ena(vcc),
	.q(\baud_rate_counter[7]~q ),
	.prn(vcc));
defparam \baud_rate_counter[7] .is_wysiwyg = "true";
defparam \baud_rate_counter[7] .power_up = "low";

cyclone10lp_lcell_comb \Equal0~1 (
	.dataa(\baud_rate_counter[4]~q ),
	.datab(\baud_rate_counter[5]~q ),
	.datac(\baud_rate_counter[6]~q ),
	.datad(\baud_rate_counter[7]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'h7FFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \baud_rate_counter[8]~25 (
	.dataa(\baud_rate_counter[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\baud_rate_counter[7]~24 ),
	.combout(\baud_rate_counter[8]~25_combout ),
	.cout());
defparam \baud_rate_counter[8]~25 .lut_mask = 16'h5A5A;
defparam \baud_rate_counter[8]~25 .sum_lutc_input = "cin";

dffeas \baud_rate_counter[8] (
	.clk(clk),
	.d(\baud_rate_counter[8]~25_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always4~0_combout ),
	.ena(vcc),
	.q(\baud_rate_counter[8]~q ),
	.prn(vcc));
defparam \baud_rate_counter[8] .is_wysiwyg = "true";
defparam \baud_rate_counter[8] .power_up = "low";

cyclone10lp_lcell_comb \always4~0 (
	.dataa(\do_load_shifter~q ),
	.datab(\Equal0~0_combout ),
	.datac(\Equal0~1_combout ),
	.datad(\baud_rate_counter[8]~q ),
	.cin(gnd),
	.combout(\always4~0_combout ),
	.cout());
defparam \always4~0 .lut_mask = 16'hFEFF;
defparam \always4~0 .sum_lutc_input = "datac";

dffeas \baud_rate_counter[0] (
	.clk(clk),
	.d(\baud_rate_counter[0]~9_combout ),
	.asdata(GND_port),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always4~0_combout ),
	.ena(vcc),
	.q(\baud_rate_counter[0]~q ),
	.prn(vcc));
defparam \baud_rate_counter[0] .is_wysiwyg = "true";
defparam \baud_rate_counter[0] .power_up = "low";

cyclone10lp_lcell_comb \Equal0~0 (
	.dataa(\baud_rate_counter[0]~q ),
	.datab(\baud_rate_counter[1]~q ),
	.datac(\baud_rate_counter[2]~q ),
	.datad(\baud_rate_counter[3]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'h7FFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal0~2 (
	.dataa(\Equal0~0_combout ),
	.datab(\Equal0~1_combout ),
	.datac(gnd),
	.datad(\baud_rate_counter[8]~q ),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
defparam \Equal0~2 .lut_mask = 16'hEEFF;
defparam \Equal0~2 .sum_lutc_input = "datac";

dffeas baud_clk_en(
	.clk(clk),
	.d(\Equal0~2_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_clk_en~q ),
	.prn(vcc));
defparam baud_clk_en.is_wysiwyg = "true";
defparam baud_clk_en.power_up = "low";

cyclone10lp_lcell_comb \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[9]~3 (
	.dataa(\do_load_shifter~q ),
	.datab(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[9]~q ),
	.datac(gnd),
	.datad(\baud_clk_en~q ),
	.cin(gnd),
	.combout(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[9]~3_combout ),
	.cout());
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[9]~3 .lut_mask = 16'hEEFF;
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[9]~3 .sum_lutc_input = "datac";

dffeas \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[9] (
	.clk(clk),
	.d(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[9]~3_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[9]~q ),
	.prn(vcc));
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[9] .is_wysiwyg = "true";
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[9] .power_up = "low";

cyclone10lp_lcell_comb \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[8]~4 (
	.dataa(tx_data_7),
	.datab(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[9]~q ),
	.datac(gnd),
	.datad(\do_load_shifter~q ),
	.cin(gnd),
	.combout(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[8]~4_combout ),
	.cout());
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[8]~4 .lut_mask = 16'hAACC;
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[8]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[4]~1 (
	.dataa(\do_load_shifter~q ),
	.datab(\WideOr0~combout ),
	.datac(\baud_clk_en~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[4]~1_combout ),
	.cout());
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[4]~1 .lut_mask = 16'hFEFE;
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[4]~1 .sum_lutc_input = "datac";

dffeas \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[8] (
	.clk(clk),
	.d(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[8]~4_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[4]~1_combout ),
	.q(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[8]~q ),
	.prn(vcc));
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[8] .is_wysiwyg = "true";
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[8] .power_up = "low";

cyclone10lp_lcell_comb \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[7]~5 (
	.dataa(tx_data_6),
	.datab(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[8]~q ),
	.datac(gnd),
	.datad(\do_load_shifter~q ),
	.cin(gnd),
	.combout(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[7]~5_combout ),
	.cout());
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[7]~5 .lut_mask = 16'hAACC;
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[7]~5 .sum_lutc_input = "datac";

dffeas \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[7] (
	.clk(clk),
	.d(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[7]~5_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[4]~1_combout ),
	.q(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[7]~q ),
	.prn(vcc));
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[7] .is_wysiwyg = "true";
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[7] .power_up = "low";

cyclone10lp_lcell_comb \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[6]~6 (
	.dataa(tx_data_5),
	.datab(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[7]~q ),
	.datac(gnd),
	.datad(\do_load_shifter~q ),
	.cin(gnd),
	.combout(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[6]~6_combout ),
	.cout());
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[6]~6 .lut_mask = 16'hAACC;
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[6]~6 .sum_lutc_input = "datac";

dffeas \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[6] (
	.clk(clk),
	.d(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[6]~6_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[4]~1_combout ),
	.q(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[6]~q ),
	.prn(vcc));
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[6] .is_wysiwyg = "true";
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[6] .power_up = "low";

cyclone10lp_lcell_comb \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[5]~7 (
	.dataa(tx_data_4),
	.datab(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[6]~q ),
	.datac(gnd),
	.datad(\do_load_shifter~q ),
	.cin(gnd),
	.combout(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[5]~7_combout ),
	.cout());
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[5]~7 .lut_mask = 16'hAACC;
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[5]~7 .sum_lutc_input = "datac";

dffeas \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[5] (
	.clk(clk),
	.d(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[5]~7_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[4]~1_combout ),
	.q(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[5]~q ),
	.prn(vcc));
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[5] .is_wysiwyg = "true";
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[5] .power_up = "low";

cyclone10lp_lcell_comb \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[4]~8 (
	.dataa(tx_data_3),
	.datab(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[5]~q ),
	.datac(gnd),
	.datad(\do_load_shifter~q ),
	.cin(gnd),
	.combout(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[4]~8_combout ),
	.cout());
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[4]~8 .lut_mask = 16'hAACC;
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[4]~8 .sum_lutc_input = "datac";

dffeas \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[4] (
	.clk(clk),
	.d(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[4]~8_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[4]~1_combout ),
	.q(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[4]~q ),
	.prn(vcc));
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[4] .is_wysiwyg = "true";
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[4] .power_up = "low";

cyclone10lp_lcell_comb \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[3]~9 (
	.dataa(tx_data_2),
	.datab(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[4]~q ),
	.datac(gnd),
	.datad(\do_load_shifter~q ),
	.cin(gnd),
	.combout(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[3]~9_combout ),
	.cout());
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[3]~9 .lut_mask = 16'hAACC;
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[3]~9 .sum_lutc_input = "datac";

dffeas \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[3] (
	.clk(clk),
	.d(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[3]~9_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[4]~1_combout ),
	.q(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[3]~q ),
	.prn(vcc));
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[3] .is_wysiwyg = "true";
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[3] .power_up = "low";

cyclone10lp_lcell_comb \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[2]~10 (
	.dataa(tx_data_1),
	.datab(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[3]~q ),
	.datac(gnd),
	.datad(\do_load_shifter~q ),
	.cin(gnd),
	.combout(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[2]~10_combout ),
	.cout());
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[2]~10 .lut_mask = 16'hAACC;
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[2]~10 .sum_lutc_input = "datac";

dffeas \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[2] (
	.clk(clk),
	.d(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[2]~10_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[4]~1_combout ),
	.q(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[2]~q ),
	.prn(vcc));
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[2] .is_wysiwyg = "true";
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[2] .power_up = "low";

cyclone10lp_lcell_comb \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[1]~11 (
	.dataa(tx_data_0),
	.datab(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[2]~q ),
	.datac(gnd),
	.datad(\do_load_shifter~q ),
	.cin(gnd),
	.combout(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[1]~11_combout ),
	.cout());
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[1]~11 .lut_mask = 16'hAACC;
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[1]~11 .sum_lutc_input = "datac";

dffeas \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[1] (
	.clk(clk),
	.d(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[1]~11_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[4]~1_combout ),
	.q(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[1]~q ),
	.prn(vcc));
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[1] .is_wysiwyg = "true";
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[1] .power_up = "low";

cyclone10lp_lcell_comb \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[0]~0 (
	.dataa(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[1]~q ),
	.datab(\baud_clk_en~q ),
	.datac(gnd),
	.datad(\do_load_shifter~q ),
	.cin(gnd),
	.combout(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[0]~0_combout ),
	.cout());
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[0]~0 .lut_mask = 16'hEEFF;
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[0]~2 (
	.dataa(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[0]~0_combout ),
	.datab(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[0]~q ),
	.datac(gnd),
	.datad(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[4]~1_combout ),
	.cin(gnd),
	.combout(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[0]~2_combout ),
	.cout());
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[0]~2 .lut_mask = 16'hEEFF;
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[0]~2 .sum_lutc_input = "datac";

dffeas \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[0] (
	.clk(clk),
	.d(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_in[0]~2_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[0]~q ),
	.prn(vcc));
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[0] .is_wysiwyg = "true";
defparam \unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[0] .power_up = "low";

cyclone10lp_lcell_comb \pre_txd~2 (
	.dataa(\pre_txd~0_combout ),
	.datab(\pre_txd~1_combout ),
	.datac(\pre_txd~q ),
	.datad(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[1]~q ),
	.cin(gnd),
	.combout(\pre_txd~2_combout ),
	.cout());
defparam \pre_txd~2 .lut_mask = 16'hEFFF;
defparam \pre_txd~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_txd~3 (
	.dataa(\unxshiftxtx_shift_register_contentsxtx_shift_reg_outxx5_out[0]~q ),
	.datab(\pre_txd~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_txd~3_combout ),
	.cout());
defparam \pre_txd~3 .lut_mask = 16'h7777;
defparam \pre_txd~3 .sum_lutc_input = "datac";

dffeas pre_txd(
	.clk(clk),
	.d(\pre_txd~3_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pre_txd~q ),
	.prn(vcc));
defparam pre_txd.is_wysiwyg = "true";
defparam pre_txd.power_up = "low";

cyclone10lp_lcell_comb \txd~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\pre_txd~q ),
	.datad(control_reg_9),
	.cin(gnd),
	.combout(\txd~0_combout ),
	.cout());
defparam \txd~0 .lut_mask = 16'hFFF0;
defparam \txd~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \tx_ready~0 (
	.dataa(\do_load_shifter~q ),
	.datab(end_begintransfer),
	.datac(tx_wr_strobe_onset1),
	.datad(tx_ready1),
	.cin(gnd),
	.combout(\tx_ready~0_combout ),
	.cout());
defparam \tx_ready~0 .lut_mask = 16'hFFF7;
defparam \tx_ready~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \tx_overrun~0 (
	.dataa(tx_wr_strobe_onset),
	.datab(tx_ready1),
	.datac(Equal2),
	.datad(end_begintransfer),
	.cin(gnd),
	.combout(\tx_overrun~0_combout ),
	.cout());
defparam \tx_overrun~0 .lut_mask = 16'hFEFF;
defparam \tx_overrun~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \tx_overrun~1 (
	.dataa(tx_overrun1),
	.datab(\tx_overrun~0_combout ),
	.datac(gnd),
	.datad(status_wr_strobe),
	.cin(gnd),
	.combout(\tx_overrun~1_combout ),
	.cout());
defparam \tx_overrun~1 .lut_mask = 16'hEEFF;
defparam \tx_overrun~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \tx_shift_empty~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\WideOr0~combout ),
	.datad(tx_ready1),
	.cin(gnd),
	.combout(\tx_shift_empty~0_combout ),
	.cout());
defparam \tx_shift_empty~0 .lut_mask = 16'hFFF0;
defparam \tx_shift_empty~0 .sum_lutc_input = "datac";

endmodule
